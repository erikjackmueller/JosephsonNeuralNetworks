* lib of neuron relevant circuits

.SUBCKT Neuron-Soma	0	1	6
* inductances
L0	0	1	3.34pH
L1	2	3	0.51pH
L2	3	4	1.09pH
L3	4	5	4.41pH
L4	5	6	2.21pH

* junctions
B0	1	2	jsoma
B1	4	0	jsoma	
B2	5	0	jsoma ic=250uA

* sources
IB0	0	3	277uA
IB1	0	5	175uA

.model jsoma jj(rtype=0, icrit=225.000uA cap=1.2PF RN=0.925)
.ends Neuron-Soma

.SUBCKT Delay-JTL	0	1	5
* inductances
L0	1	2	2.127pH
L1	2	3	2.080pH
L2	3	4	2.080pH
L3	4	5	2.127pH

* junctions
B0	2	0	jdelay 
B1	4	0	jdelay 

* sources
IB0	0	3	250uA

.model jdelay jj(rtype=0, icrit=250.000uA cap=1.2PF RN=0.877)
.ends Delay-JTL


.SUBCKT JJ-Soma	0	1	3
* inductances
L0	1	2	1.0pH
L1	2	3 	1.0pH

* junctions
B0	2	0	jj1

* sources
IB0 	0	2 	175uA

.model jj1 jj(rtype=0, icrit=250.000uA cap=4PF RN=0.877)
.ends JJ-Soma

.SUBCKT R-Synapse-exc	0	1	2
* inductances
R1	1	0	1
RSCALE	1	2	1
.ends R-Synapse-exc

.SUBCKT R-Synapse-inh	0	1	5
* inductances
L0	1	2	1.0pH
L1	3	4	1.0pH
R1	4	0	1.0 
RSCALE	4	5	1.0
* this should function as the same scaling output as in the exc case

* junctions
B0	2	3	jsyn ic=200uA
B1	3	0	jsyn ic=1000uA

.model jsyn jj(rtype=0, icrit=250.000uA cap=1.2PF RN=0.877)
.ends R-Synapse-inh


.SUBCKT 2-Split	0	1	6	8
* inductances
L1	1	2	1.183pH
L2	2	3	1.420pH
L3	3	4	0.509pH
L4	4	5	1.679pH
L5	5	6	1.900pH
L6	4	7	1.634pH
L7	7	8	1.897pH

* junctions
B1	2	0	jsplit ic=325uA
B2	5	0	jsplit 
B3	7	0	jsplit 

* sources
IB	0	3	570uA

.model jsplit jj(rtype=0, icrit=250.000uA cap=1.2PF RN=0.877)
.ends 2-Split

.SUBCKT 3-Split	0	1	6	8	10
* inductances
L1	1	2	1.183pH
L2	2	3	1.420pH
L3	3	4	0.509pH
L4	4	5	1.650pH
L5	5	6	1.900pH
L6	4	7	1.650pH
L7	7	8	1.900pH
*-------------------------------
L8	4	9	1.650pH
L9	9	10	1.900pH

* junctions
B1	2	0	jsplit ic=325uA
B2	5	0	jsplit 
B3	7	0	jsplit 
*-------------------------------
B4	9	0	jsplit

* sources
IB	0	3	855uA
* 570*1.5

.model jsplit jj(rtype=0, icrit=250.000uA cap=1.2PF RN=0.877)
.ends 3-Split







* Josim Circuit automatically assembled using build_circuit on 2025-07-01 14:05:26.897988 
 
.SUBCKT exc-neuron	0	1	2	3	4	5	6	7	8	9	10	11	
 
X0	Neuron-Soma	0	1	soma-split	
X1	2-Split	0	soma-split	2_syn	3_syn	4_syn	5_syn	6_syn	7_syn	8_syn	9_syn	10_syn	11_syn	
X2	R-Synapse-exc	0	2_syn	2	
X3	R-Synapse-exc	0	3_syn	3	
X4	R-Synapse-exc	0	4_syn	4	
X5	R-Synapse-exc	0	5_syn	5	
X6	R-Synapse-exc	0	6_syn	6	
X7	R-Synapse-exc	0	7_syn	7	
X8	R-Synapse-exc	0	8_syn	8	
X9	R-Synapse-exc	0	9_syn	9	
X10	R-Synapse-exc	0	10_syn	10	
X11	R-Synapse-exc	0	11_syn	11	
.ends exc-neuron

.SUBCKT R-Synapse-exc	0	1	2
* inductances
R1	1	0	1
RSCALE	1	2	1
.ends R-Synapse-exc

.SUBCKT 2-Split	0	1	6	8	10	12	14	16	18	20	22	24
* inductances
L1	1	2	1.183pH
L2	2	3	1.420pH
L3	3	4	0.509pH
L4	4	5	1.679pH
L5	5	6	1.900pH
L6	4	7	1.634pH
L7	7	8	1.897pH
L8	4	9	1.65pH
L9	9	10	1.9pH
L10	4	11	1.65pH
L11	11	12	1.9pH
L12	4	13	1.65pH
L13	13	14	1.9pH
L14	4	15	1.65pH
L15	15	16	1.9pH
L16	4	17	1.65pH
L17	17	18	1.9pH
L18	4	19	1.65pH
L19	19	20	1.9pH
L20	4	21	1.65pH
L21	21	22	1.9pH
L22	4	23	1.65pH
L23	23	24	1.9pH

* junctions
B1	2	0	jsplit ic=325uA
B2	5	0	jsplit 
B3	7	0	jsplit 
B4	9	0	jsplit
B5	11	0	jsplit
B6	13	0	jsplit
B7	15	0	jsplit
B8	17	0	jsplit
B9	19	0	jsplit
B10	21	0	jsplit
B11	23	0	jsplit

* sources
IB	0	3	2850.0uA
.model jsplit jj(rtype=0, icrit=250.000uA cap=1.2PF RN=0.877)
.ends 2-Split

.SUBCKT Neuron-Soma	0	1	6
* inductances
L0	0	1	3.34pH
L1	2	3	0.51pH
L2	3	4	1.09pH
L3	4	5	4.41pH
L4	5	6	2.21pH

* junctions
B0	1	2	jsoma
B1	4	0	jsoma	
B2	5	0	jsoma ic=250uA

* sources
IB0	0	3	277uA
IB1	0	5	175uA

.model jsoma jj(rtype=0, icrit=225.000uA cap=1.2PF RN=0.925)
.ends Neuron-Soma


* main circuit
IIN0 0 1 pwl(0 0 0.764p 0 0.765p 10000.0u 0.766p 0 10.283p 0 10.284p 10000.0u 10.285p 0 11.651p 0 11.652p 10000.0u 11.653p 0 29.837p 0 29.838p 10000.0u 29.839p 0 39.407p 0 39.408p 10000.0u 39.409p 0 42.014p 0 42.015p 10000.0u 42.016p 0 71.129p 0 71.13p 10000.0u 71.131p 0 82.904p 0 82.905p 10000.0u 82.906p 0 83.066p 0 83.067p 10000.0u 83.068p 0 83.273p 0 83.274p 10000.0u 83.275p 0 89.555p 0 89.556p 10000.0u 89.557p 0 95.261p 0 95.262p 10000.0u 95.263p 0 129.734p 0 129.735p 10000.0u 129.736p 0 138.755p 0 138.756p 10000.0u 138.757p 0 142.484p 0 142.485p 10000.0u 142.486p 0 144.377p 0 144.378p 10000.0u 144.379p 0 149.231p 0 149.232p 10000.0u 149.233p 0 150.302p 0 150.303p 10000.0u 150.304p 0 160.022p 0 160.023p 10000.0u 160.024p 0 180.296p 0 180.297p 10000.0u 180.298p 0 181.199p 0 181.2p 10000.0u 181.201p 0 183.974p 0 183.975p 10000.0u 183.976p 0 187.838p 0 187.839p 10000.0u 187.84p 0 188.273p 0 188.274p 10000.0u 188.275p 0 197.285p 0 197.286p 10000.0u 197.287p 0 205.208p 0 205.209p 10000.0u 205.21p 0 220.973p 0 220.974p 10000.0u 220.975p 0 224.807p 0 224.808p 10000.0u 224.809p 0 226.007p 0 226.008p 10000.0u 226.009p 0 232.277p 0 232.278p 10000.0u 232.279p 0 240.317p 0 240.318p 10000.0u 240.319p 0 250.226p 0 250.227p 10000.0u 250.228p 0 253.7p 0 253.701p 10000.0u 253.702p 0 267.551p 0 267.552p 10000.0u 267.553p 0 268.529p 0 268.53p 10000.0u 268.531p 0 270.776p 0 270.777p 10000.0u 270.778p 0 287.273p 0 287.274p 10000.0u 287.275p 0 295.106p 0 295.107p 10000.0u 295.108p 0 298.283p 0 298.284p 10000.0u 298.285p 0 300.911p 0 300.912p 10000.0u 300.913p 0 327.044p 0 327.045p 10000.0u 327.046p 0 370.127p 0 370.128p 10000.0u 370.129p 0 378.41p 0 378.411p 10000.0u 378.412p 0 386.549p 0 386.55p 10000.0u 386.551p 0 389.318p 0 389.319p 10000.0u 389.32p 0 403.175p 0 403.176p 10000.0u 403.177p 0 416.519p 0 416.52p 10000.0u 416.521p 0 433.19p 0 433.191p 10000.0u 433.192p 0 449.243p 0 449.244p 10000.0u 449.245p 0 451.655p 0 451.656p 10000.0u 451.657p 0 456.491p 0 456.492p 10000.0u 456.493p 0 459.365p 0 459.366p 10000.0u 459.367p 0 460.961p 0 460.962p 10000.0u 460.963p 0 461.306p 0 461.307p 10000.0u 461.308p 0 486.845p 0 486.846p 10000.0u 486.847p 0 508.886p 0 508.887p 10000.0u 508.888p 0 519.536p 0 519.537p 10000.0u 519.538p 0 524.993p 0 524.994p 10000.0u 524.995p 0 533.051p 0 533.052p 10000.0u 533.053p 0 569.861p 0 569.862p 10000.0u 569.863p 0 573.659p 0 573.66p 10000.0u 573.661p 0 580.205p 0 580.206p 10000.0u 580.207p 0 593.186p 0 593.187p 10000.0u 593.188p 0 596.012p 0 596.013p 10000.0u 596.014p 0 602.06p 0 602.061p 10000.0u 602.062p 0 615.602p 0 615.603p 10000.0u 615.604p 0 621.611p 0 621.612p 10000.0u 621.613p 0 627.311p 0 627.312p 10000.0u 627.313p 0 628.028p 0 628.029p 10000.0u 628.03p 0 628.79p 0 628.791p 10000.0u 628.792p 0 636.134p 0 636.135p 10000.0u 636.136p 0 642.641p 0 642.642p 10000.0u 642.643p 0 650.474p 0 650.475p 10000.0u 650.476p 0 659.222p 0 659.223p 10000.0u 659.224p 0 668.618p 0 668.619p 10000.0u 668.62p 0 674.333p 0 674.334p 10000.0u 674.335p 0 676.448p 0 676.449p 10000.0u 676.45p 0 691.493p 0 691.494p 10000.0u 691.495p 0 694.664p 0 694.665p 10000.0u 694.666p 0 739.646p 0 739.647p 10000.0u 739.648p 0 745.295p 0 745.296p 10000.0u 745.297p 0 755.714p 0 755.715p 10000.0u 755.716p 0 764.615p 0 764.616p 10000.0u 764.617p 0 776.78p 0 776.781p 10000.0u 776.782p 0 777.791p 0 777.792p 10000.0u 777.793p 0 788.594p 0 788.595p 10000.0u 788.596p 0 789.308p 0 789.309p 10000.0u 789.31p 0 791.018p 0 791.019p 10000.0u 791.02p 0 792.59p 0 792.591p 10000.0u 792.592p 0 808.79p 0 808.791p 10000.0u 808.792p 0 820.316p 0 820.317p 10000.0u 820.318p 0 823.214p 0 823.215p 10000.0u 823.216p 0 882.101p 0 882.102p 10000.0u 882.103p 0 899.675p 0 899.676p 10000.0u 899.677p 0 917.309p 0 917.31p 10000.0u 917.311p 0 933.446p 0 933.447p 10000.0u 933.448p 0 948.866p 0 948.867p 10000.0u 948.868p 0 956.849p 0 956.85p 10000.0u 956.851p 0 960.419p 0 960.42p 10000.0u 960.421p 0 960.581p 0 960.582p 10000.0u 960.583p 0 963.35p 0 963.351p 10000.0u 963.352p 0 985.253p 0 985.254p 10000.0u 985.255p 0)
IIN1 0 2 pwl(0 0 51.323p 0 51.324p 10000.0u 51.325p 0 60.104p 0 60.105p 10000.0u 60.106p 0 76.259p 0 76.26p 10000.0u 76.261p 0 83.096p 0 83.097p 10000.0u 83.098p 0 88.265p 0 88.266p 10000.0u 88.267p 0 89.249p 0 89.25p 10000.0u 89.251p 0 104.909p 0 104.91p 10000.0u 104.911p 0 107.261p 0 107.262p 10000.0u 107.263p 0 109.271p 0 109.272p 10000.0u 109.273p 0 111.524p 0 111.525p 10000.0u 111.526p 0 123.128p 0 123.129p 10000.0u 123.13p 0 139.151p 0 139.152p 10000.0u 139.153p 0 139.52p 0 139.521p 10000.0u 139.522p 0 150.521p 0 150.522p 10000.0u 150.523p 0 155.111p 0 155.112p 10000.0u 155.113p 0 165.467p 0 165.468p 10000.0u 165.469p 0 180.368p 0 180.369p 10000.0u 180.37p 0 183.959p 0 183.96p 10000.0u 183.961p 0 207.311p 0 207.312p 10000.0u 207.313p 0 208.841p 0 208.842p 10000.0u 208.843p 0 213.371p 0 213.372p 10000.0u 213.373p 0 226.793p 0 226.794p 10000.0u 226.795p 0 236.336p 0 236.337p 10000.0u 236.338p 0 237.698p 0 237.699p 10000.0u 237.7p 0 251.141p 0 251.142p 10000.0u 251.143p 0 254.159p 0 254.16p 10000.0u 254.161p 0 259.13p 0 259.131p 10000.0u 259.132p 0 259.193p 0 259.194p 10000.0u 259.195p 0 265.673p 0 265.674p 10000.0u 265.675p 0 304.58p 0 304.581p 10000.0u 304.582p 0 307.253p 0 307.254p 10000.0u 307.255p 0 313.814p 0 313.815p 10000.0u 313.816p 0 314.378p 0 314.379p 10000.0u 314.38p 0 328.016p 0 328.017p 10000.0u 328.018p 0 329.738p 0 329.739p 10000.0u 329.74p 0 330.857p 0 330.858p 10000.0u 330.859p 0 361.556p 0 361.557p 10000.0u 361.558p 0 370.433p 0 370.434p 10000.0u 370.435p 0 376.085p 0 376.086p 10000.0u 376.087p 0 387.383p 0 387.384p 10000.0u 387.385p 0 392.969p 0 392.97p 10000.0u 392.971p 0 403.376p 0 403.377p 10000.0u 403.378p 0 418.352p 0 418.353p 10000.0u 418.354p 0 427.451p 0 427.452p 10000.0u 427.453p 0 438.476p 0 438.477p 10000.0u 438.478p 0 459.944p 0 459.945p 10000.0u 459.946p 0 475.586p 0 475.587p 10000.0u 475.588p 0 483.194p 0 483.195p 10000.0u 483.196p 0 485.003p 0 485.004p 10000.0u 485.005p 0 514.781p 0 514.782p 10000.0u 514.783p 0 521.411p 0 521.412p 10000.0u 521.413p 0 531.818p 0 531.819p 10000.0u 531.82p 0 532.97p 0 532.971p 10000.0u 532.972p 0 539.45p 0 539.451p 10000.0u 539.452p 0 540.098p 0 540.099p 10000.0u 540.1p 0 563.9p 0 563.901p 10000.0u 563.902p 0 571.874p 0 571.875p 10000.0u 571.876p 0 584.393p 0 584.394p 10000.0u 584.395p 0 605.558p 0 605.559p 10000.0u 605.56p 0 609.56p 0 609.561p 10000.0u 609.562p 0 616.511p 0 616.512p 10000.0u 616.513p 0 617.045p 0 617.046p 10000.0u 617.047p 0 624.434p 0 624.435p 10000.0u 624.436p 0 625.973p 0 625.974p 10000.0u 625.975p 0 638.555p 0 638.556p 10000.0u 638.557p 0 665.837p 0 665.838p 10000.0u 665.839p 0 671.987p 0 671.988p 10000.0u 671.989p 0 672.716p 0 672.717p 10000.0u 672.718p 0 673.829p 0 673.83p 10000.0u 673.831p 0 686.426p 0 686.427p 10000.0u 686.428p 0 689.855p 0 689.856p 10000.0u 689.857p 0 697.451p 0 697.452p 10000.0u 697.453p 0 722.153p 0 722.154p 10000.0u 722.155p 0 729.962p 0 729.963p 10000.0u 729.964p 0 730.979p 0 730.98p 10000.0u 730.981p 0 741.038p 0 741.039p 10000.0u 741.04p 0 745.886p 0 745.887p 10000.0u 745.888p 0 785.528p 0 785.529p 10000.0u 785.53p 0 815.51p 0 815.511p 10000.0u 815.512p 0 839.627p 0 839.628p 10000.0u 839.629p 0 843.371p 0 843.372p 10000.0u 843.373p 0 870.143p 0 870.144p 10000.0u 870.145p 0 871.241p 0 871.242p 10000.0u 871.243p 0 892.796p 0 892.797p 10000.0u 892.798p 0 896.288p 0 896.289p 10000.0u 896.29p 0 896.849p 0 896.85p 10000.0u 896.851p 0 903.719p 0 903.72p 10000.0u 903.721p 0 919.106p 0 919.107p 10000.0u 919.108p 0 936.404p 0 936.405p 10000.0u 936.406p 0 938.033p 0 938.034p 10000.0u 938.035p 0 938.702p 0 938.703p 10000.0u 938.704p 0 939.674p 0 939.675p 10000.0u 939.676p 0 943.97p 0 943.971p 10000.0u 943.972p 0 955.163p 0 955.164p 10000.0u 955.165p 0 969.686p 0 969.687p 10000.0u 969.688p 0 990.047p 0 990.048p 10000.0u 990.049p 0 994.655p 0 994.656p 10000.0u 994.657p 0)
IIN2 0 3 pwl(0 0 1.904p 0 1.905p 10000.0u 1.906p 0 19.559p 0 19.56p 10000.0u 19.561p 0 26.798p 0 26.799p 10000.0u 26.8p 0 46.4p 0 46.401p 10000.0u 46.402p 0 47.951p 0 47.952p 10000.0u 47.953p 0 52.895p 0 52.896p 10000.0u 52.897p 0 56.672p 0 56.673p 10000.0u 56.674p 0 110.042p 0 110.043p 10000.0u 110.044p 0 126.785p 0 126.786p 10000.0u 126.787p 0 136.031p 0 136.032p 10000.0u 136.033p 0 143.633p 0 143.634p 10000.0u 143.635p 0 149.45p 0 149.451p 10000.0u 149.452p 0 182.18p 0 182.181p 10000.0u 182.182p 0 182.414p 0 182.415p 10000.0u 182.416p 0 187.055p 0 187.056p 10000.0u 187.057p 0 190.331p 0 190.332p 10000.0u 190.333p 0 194.117p 0 194.118p 10000.0u 194.119p 0 202.769p 0 202.77p 10000.0u 202.771p 0 208.301p 0 208.302p 10000.0u 208.303p 0 209.498p 0 209.499p 10000.0u 209.5p 0 227.186p 0 227.187p 10000.0u 227.188p 0 232.715p 0 232.716p 10000.0u 232.717p 0 239.315p 0 239.316p 10000.0u 239.317p 0 247.892p 0 247.893p 10000.0u 247.894p 0 248.954p 0 248.955p 10000.0u 248.956p 0 253.025p 0 253.026p 10000.0u 253.027p 0 255.509p 0 255.51p 10000.0u 255.511p 0 257.501p 0 257.502p 10000.0u 257.503p 0 258.212p 0 258.213p 10000.0u 258.214p 0 267.983p 0 267.984p 10000.0u 267.985p 0 282.578p 0 282.579p 10000.0u 282.58p 0 286.961p 0 286.962p 10000.0u 286.963p 0 291.239p 0 291.24p 10000.0u 291.241p 0 296.348p 0 296.349p 10000.0u 296.35p 0 302.465p 0 302.466p 10000.0u 302.467p 0 306.347p 0 306.348p 10000.0u 306.349p 0 334.022p 0 334.023p 10000.0u 334.024p 0 344.192p 0 344.193p 10000.0u 344.194p 0 373.319p 0 373.32p 10000.0u 373.321p 0 384.59p 0 384.591p 10000.0u 384.592p 0 394.913p 0 394.914p 10000.0u 394.915p 0 409.265p 0 409.266p 10000.0u 409.267p 0 409.565p 0 409.566p 10000.0u 409.567p 0 410.96p 0 410.961p 10000.0u 410.962p 0 440.045p 0 440.046p 10000.0u 440.047p 0 452.474p 0 452.475p 10000.0u 452.476p 0 452.921p 0 452.922p 10000.0u 452.923p 0 454.697p 0 454.698p 10000.0u 454.699p 0 467.714p 0 467.715p 10000.0u 467.716p 0 478.499p 0 478.5p 10000.0u 478.501p 0 488.498p 0 488.499p 10000.0u 488.5p 0 491.258p 0 491.259p 10000.0u 491.26p 0 499.694p 0 499.695p 10000.0u 499.696p 0 502.736p 0 502.737p 10000.0u 502.738p 0 505.691p 0 505.692p 10000.0u 505.693p 0 515.819p 0 515.82p 10000.0u 515.821p 0 531.311p 0 531.312p 10000.0u 531.313p 0 533.753p 0 533.754p 10000.0u 533.755p 0 537.155p 0 537.156p 10000.0u 537.157p 0 564.761p 0 564.762p 10000.0u 564.763p 0 565.937p 0 565.938p 10000.0u 565.939p 0 573.77p 0 573.771p 10000.0u 573.772p 0 574.271p 0 574.272p 10000.0u 574.273p 0 580.229p 0 580.23p 10000.0u 580.231p 0 590.699p 0 590.7p 10000.0u 590.701p 0 595.679p 0 595.68p 10000.0u 595.681p 0 633.365p 0 633.366p 10000.0u 633.367p 0 640.007p 0 640.008p 10000.0u 640.009p 0 643.823p 0 643.824p 10000.0u 643.825p 0 644.519p 0 644.52p 10000.0u 644.521p 0 650.591p 0 650.592p 10000.0u 650.593p 0 653.822p 0 653.823p 10000.0u 653.824p 0 656.582p 0 656.583p 10000.0u 656.584p 0 662.474p 0 662.475p 10000.0u 662.476p 0 672.023p 0 672.024p 10000.0u 672.025p 0 674.105p 0 674.106p 10000.0u 674.107p 0 701.252p 0 701.253p 10000.0u 701.254p 0 704.642p 0 704.643p 10000.0u 704.644p 0 716.582p 0 716.583p 10000.0u 716.584p 0 726.653p 0 726.654p 10000.0u 726.655p 0 735.878p 0 735.879p 10000.0u 735.88p 0 775.154p 0 775.155p 10000.0u 775.156p 0 794.189p 0 794.19p 10000.0u 794.191p 0 799.121p 0 799.122p 10000.0u 799.123p 0 801.296p 0 801.297p 10000.0u 801.298p 0 812.354p 0 812.355p 10000.0u 812.356p 0 812.633p 0 812.634p 10000.0u 812.635p 0 828.494p 0 828.495p 10000.0u 828.496p 0 848.831p 0 848.832p 10000.0u 848.833p 0 852.953p 0 852.954p 10000.0u 852.955p 0 855.026p 0 855.027p 10000.0u 855.028p 0 855.935p 0 855.936p 10000.0u 855.937p 0 867.368p 0 867.369p 10000.0u 867.37p 0 960.782p 0 960.783p 10000.0u 960.784p 0 982.571p 0 982.572p 10000.0u 982.573p 0 986.597p 0 986.598p 10000.0u 986.599p 0)
IIN3 0 4 pwl(0 0 21.644p 0 21.645p 10000.0u 21.646p 0 29.777p 0 29.778p 10000.0u 29.779p 0 50.183p 0 50.184p 10000.0u 50.185p 0 53.132p 0 53.133p 10000.0u 53.134p 0 55.481p 0 55.482p 10000.0u 55.483p 0 76.034p 0 76.035p 10000.0u 76.036p 0 87.071p 0 87.072p 10000.0u 87.073p 0 98.372p 0 98.373p 10000.0u 98.374p 0 99.926p 0 99.927p 10000.0u 99.928p 0 100.673p 0 100.674p 10000.0u 100.675p 0 115.937p 0 115.938p 10000.0u 115.939p 0 127.817p 0 127.818p 10000.0u 127.819p 0 137.384p 0 137.385p 10000.0u 137.386p 0 151.823p 0 151.824p 10000.0u 151.825p 0 158.255p 0 158.256p 10000.0u 158.257p 0 163.085p 0 163.086p 10000.0u 163.087p 0 164.804p 0 164.805p 10000.0u 164.806p 0 165.155p 0 165.156p 10000.0u 165.157p 0 166.628p 0 166.629p 10000.0u 166.63p 0 167.807p 0 167.808p 10000.0u 167.809p 0 173.348p 0 173.349p 10000.0u 173.35p 0 197.15p 0 197.151p 10000.0u 197.152p 0 202.016p 0 202.017p 10000.0u 202.018p 0 216.707p 0 216.708p 10000.0u 216.709p 0 219.851p 0 219.852p 10000.0u 219.853p 0 231.863p 0 231.864p 10000.0u 231.865p 0 255.776p 0 255.777p 10000.0u 255.778p 0 261.323p 0 261.324p 10000.0u 261.325p 0 262.691p 0 262.692p 10000.0u 262.693p 0 272.369p 0 272.37p 10000.0u 272.371p 0 275.822p 0 275.823p 10000.0u 275.824p 0 291.029p 0 291.03p 10000.0u 291.031p 0 302.696p 0 302.697p 10000.0u 302.698p 0 309.617p 0 309.618p 10000.0u 309.619p 0 309.776p 0 309.777p 10000.0u 309.778p 0 332.567p 0 332.568p 10000.0u 332.569p 0 333.872p 0 333.873p 10000.0u 333.874p 0 341.93p 0 341.931p 10000.0u 341.932p 0 353.513p 0 353.514p 10000.0u 353.515p 0 362.501p 0 362.502p 10000.0u 362.503p 0 363.683p 0 363.684p 10000.0u 363.685p 0 367.178p 0 367.179p 10000.0u 367.18p 0 392.24p 0 392.241p 10000.0u 392.242p 0 392.426p 0 392.427p 10000.0u 392.428p 0 398.702p 0 398.703p 10000.0u 398.704p 0 406.04p 0 406.041p 10000.0u 406.042p 0 409.682p 0 409.683p 10000.0u 409.684p 0 423.86p 0 423.861p 10000.0u 423.862p 0 425.294p 0 425.295p 10000.0u 425.296p 0 429.11p 0 429.111p 10000.0u 429.112p 0 441.854p 0 441.855p 10000.0u 441.856p 0 446.864p 0 446.865p 10000.0u 446.866p 0 450.461p 0 450.462p 10000.0u 450.463p 0 462.74p 0 462.741p 10000.0u 462.742p 0 468.938p 0 468.939p 10000.0u 468.94p 0 470.708p 0 470.709p 10000.0u 470.71p 0 483.935p 0 483.936p 10000.0u 483.937p 0 484.934p 0 484.935p 10000.0u 484.936p 0 485.639p 0 485.64p 10000.0u 485.641p 0 493.145p 0 493.146p 10000.0u 493.147p 0 504.947p 0 504.948p 10000.0u 504.949p 0 507.203p 0 507.204p 10000.0u 507.205p 0 515.186p 0 515.187p 10000.0u 515.188p 0 517.544p 0 517.545p 10000.0u 517.546p 0 521.405p 0 521.406p 10000.0u 521.407p 0 526.433p 0 526.434p 10000.0u 526.435p 0 546.512p 0 546.513p 10000.0u 546.514p 0 558.008p 0 558.009p 10000.0u 558.01p 0 565.415p 0 565.416p 10000.0u 565.417p 0 647.222p 0 647.223p 10000.0u 647.224p 0 653.261p 0 653.262p 10000.0u 653.263p 0 658.04p 0 658.041p 10000.0u 658.042p 0 668.21p 0 668.211p 10000.0u 668.212p 0 671.693p 0 671.694p 10000.0u 671.695p 0 679.436p 0 679.437p 10000.0u 679.438p 0 682.694p 0 682.695p 10000.0u 682.696p 0 683.012p 0 683.013p 10000.0u 683.014p 0 690.074p 0 690.075p 10000.0u 690.076p 0 697.253p 0 697.254p 10000.0u 697.255p 0 704.75p 0 704.751p 10000.0u 704.752p 0 713.516p 0 713.517p 10000.0u 713.518p 0 720.461p 0 720.462p 10000.0u 720.463p 0 720.71p 0 720.711p 10000.0u 720.712p 0 726.401p 0 726.402p 10000.0u 726.403p 0 750.515p 0 750.516p 10000.0u 750.517p 0 779.426p 0 779.427p 10000.0u 779.428p 0 784.13p 0 784.131p 10000.0u 784.132p 0 794.417p 0 794.418p 10000.0u 794.419p 0 804.344p 0 804.345p 10000.0u 804.346p 0 811.28p 0 811.281p 10000.0u 811.282p 0 814.592p 0 814.593p 10000.0u 814.594p 0 818.339p 0 818.34p 10000.0u 818.341p 0 833.75p 0 833.751p 10000.0u 833.752p 0 838.205p 0 838.206p 10000.0u 838.207p 0 844.46p 0 844.461p 10000.0u 844.462p 0 847.859p 0 847.86p 10000.0u 847.861p 0 851.276p 0 851.277p 10000.0u 851.278p 0 853.526p 0 853.527p 10000.0u 853.528p 0 865.643p 0 865.644p 10000.0u 865.645p 0 879.836p 0 879.837p 10000.0u 879.838p 0 901.01p 0 901.011p 10000.0u 901.012p 0 907.556p 0 907.557p 10000.0u 907.558p 0 925.493p 0 925.494p 10000.0u 925.495p 0 925.748p 0 925.749p 10000.0u 925.75p 0 934.328p 0 934.329p 10000.0u 934.33p 0 935.297p 0 935.298p 10000.0u 935.299p 0 939.584p 0 939.585p 10000.0u 939.586p 0 955.241p 0 955.242p 10000.0u 955.243p 0 956.723p 0 956.724p 10000.0u 956.725p 0 965.33p 0 965.331p 10000.0u 965.332p 0 967.655p 0 967.656p 10000.0u 967.657p 0 974.837p 0 974.838p 10000.0u 974.839p 0)
IIN4 0 5 pwl(0 0 1.817p 0 1.818p 10000.0u 1.819p 0 10.955p 0 10.956p 10000.0u 10.957p 0 16.343p 0 16.344p 10000.0u 16.345p 0 21.152p 0 21.153p 10000.0u 21.154p 0 27.2p 0 27.201p 10000.0u 27.202p 0 73.928p 0 73.929p 10000.0u 73.93p 0 74.87p 0 74.871p 10000.0u 74.872p 0 74.948p 0 74.949p 10000.0u 74.95p 0 96.809p 0 96.81p 10000.0u 96.811p 0 113.015p 0 113.016p 10000.0u 113.017p 0 115.025p 0 115.026p 10000.0u 115.027p 0 115.664p 0 115.665p 10000.0u 115.666p 0 144.698p 0 144.699p 10000.0u 144.7p 0 160.136p 0 160.137p 10000.0u 160.138p 0 160.547p 0 160.548p 10000.0u 160.549p 0 167.867p 0 167.868p 10000.0u 167.869p 0 170.135p 0 170.136p 10000.0u 170.137p 0 174.029p 0 174.03p 10000.0u 174.031p 0 183.389p 0 183.39p 10000.0u 183.391p 0 193.937p 0 193.938p 10000.0u 193.939p 0 199.688p 0 199.689p 10000.0u 199.69p 0 209.375p 0 209.376p 10000.0u 209.377p 0 228.044p 0 228.045p 10000.0u 228.046p 0 229.22p 0 229.221p 10000.0u 229.222p 0 244.256p 0 244.257p 10000.0u 244.258p 0 252.488p 0 252.489p 10000.0u 252.49p 0 270.653p 0 270.654p 10000.0u 270.655p 0 279.17p 0 279.171p 10000.0u 279.172p 0 296.888p 0 296.889p 10000.0u 296.89p 0 301.07p 0 301.071p 10000.0u 301.072p 0 303.281p 0 303.282p 10000.0u 303.283p 0 304.574p 0 304.575p 10000.0u 304.576p 0 311.333p 0 311.334p 10000.0u 311.335p 0 317.018p 0 317.019p 10000.0u 317.02p 0 327.911p 0 327.912p 10000.0u 327.913p 0 328.094p 0 328.095p 10000.0u 328.096p 0 328.187p 0 328.188p 10000.0u 328.189p 0 340.856p 0 340.857p 10000.0u 340.858p 0 352.487p 0 352.488p 10000.0u 352.489p 0 356.81p 0 356.811p 10000.0u 356.812p 0 373.841p 0 373.842p 10000.0u 373.843p 0 374.102p 0 374.103p 10000.0u 374.104p 0 418.685p 0 418.686p 10000.0u 418.687p 0 432.197p 0 432.198p 10000.0u 432.199p 0 439.292p 0 439.293p 10000.0u 439.294p 0 442.55p 0 442.551p 10000.0u 442.552p 0 451.373p 0 451.374p 10000.0u 451.375p 0 453.131p 0 453.132p 10000.0u 453.133p 0 454.928p 0 454.929p 10000.0u 454.93p 0 455.705p 0 455.706p 10000.0u 455.707p 0 458.612p 0 458.613p 10000.0u 458.614p 0 458.759p 0 458.76p 10000.0u 458.761p 0 491.411p 0 491.412p 10000.0u 491.413p 0 507.59p 0 507.591p 10000.0u 507.592p 0 512.03p 0 512.031p 10000.0u 512.032p 0 520.475p 0 520.476p 10000.0u 520.477p 0 534.266p 0 534.267p 10000.0u 534.268p 0 537.512p 0 537.513p 10000.0u 537.514p 0 538.403p 0 538.404p 10000.0u 538.405p 0 543.314p 0 543.315p 10000.0u 543.316p 0 544.754p 0 544.755p 10000.0u 544.756p 0 560.132p 0 560.133p 10000.0u 560.134p 0 566.312p 0 566.313p 10000.0u 566.314p 0 571.025p 0 571.026p 10000.0u 571.027p 0 572.123p 0 572.124p 10000.0u 572.125p 0 581.612p 0 581.613p 10000.0u 581.614p 0 582.176p 0 582.177p 10000.0u 582.178p 0 589.724p 0 589.725p 10000.0u 589.726p 0 593.081p 0 593.082p 10000.0u 593.083p 0 597.656p 0 597.657p 10000.0u 597.658p 0 617.507p 0 617.508p 10000.0u 617.509p 0 621.008p 0 621.009p 10000.0u 621.01p 0 627.761p 0 627.762p 10000.0u 627.763p 0 639.074p 0 639.075p 10000.0u 639.076p 0 650.192p 0 650.193p 10000.0u 650.194p 0 652.661p 0 652.662p 10000.0u 652.663p 0 657.722p 0 657.723p 10000.0u 657.724p 0 673.616p 0 673.617p 10000.0u 673.618p 0 681.074p 0 681.075p 10000.0u 681.076p 0 687.596p 0 687.597p 10000.0u 687.598p 0 702.713p 0 702.714p 10000.0u 702.715p 0 723.734p 0 723.735p 10000.0u 723.736p 0 726.476p 0 726.477p 10000.0u 726.478p 0 728.51p 0 728.511p 10000.0u 728.512p 0 737.123p 0 737.124p 10000.0u 737.125p 0 748.307p 0 748.308p 10000.0u 748.309p 0 748.442p 0 748.443p 10000.0u 748.444p 0 754.241p 0 754.242p 10000.0u 754.243p 0 758.537p 0 758.538p 10000.0u 758.539p 0 771.602p 0 771.603p 10000.0u 771.604p 0 778.109p 0 778.11p 10000.0u 778.111p 0 801.464p 0 801.465p 10000.0u 801.466p 0 826.856p 0 826.857p 10000.0u 826.858p 0 840.29p 0 840.291p 10000.0u 840.292p 0 846.56p 0 846.561p 10000.0u 846.562p 0 857.822p 0 857.823p 10000.0u 857.824p 0 882.431p 0 882.432p 10000.0u 882.433p 0 891.059p 0 891.06p 10000.0u 891.061p 0 898.166p 0 898.167p 10000.0u 898.168p 0 917.126p 0 917.127p 10000.0u 917.128p 0 957.545p 0 957.546p 10000.0u 957.547p 0 963.263p 0 963.264p 10000.0u 963.265p 0 975.53p 0 975.531p 10000.0u 975.532p 0 990.536p 0 990.537p 10000.0u 990.538p 0 999.608p 0 999.609p 10000.0u 999.61p 0)
IIN5 0 6 pwl(0 0 3.935p 0 3.936p 10000.0u 3.937p 0 4.49p 0 4.491p 10000.0u 4.492p 0 9.119p 0 9.12p 10000.0u 9.121p 0 14.138p 0 14.139p 10000.0u 14.14p 0 14.891p 0 14.892p 10000.0u 14.893p 0 27.158p 0 27.159p 10000.0u 27.16p 0 38.009p 0 38.01p 10000.0u 38.011p 0 41.915p 0 41.916p 10000.0u 41.917p 0 44.012p 0 44.013p 10000.0u 44.014p 0 54.71p 0 54.711p 10000.0u 54.712p 0 87.386p 0 87.387p 10000.0u 87.388p 0 91.328p 0 91.329p 10000.0u 91.33p 0 117.197p 0 117.198p 10000.0u 117.199p 0 120.563p 0 120.564p 10000.0u 120.565p 0 128.831p 0 128.832p 10000.0u 128.833p 0 129.596p 0 129.597p 10000.0u 129.598p 0 143.0p 0 143.001p 10000.0u 143.002p 0 148.892p 0 148.893p 10000.0u 148.894p 0 149.351p 0 149.352p 10000.0u 149.353p 0 165.056p 0 165.057p 10000.0u 165.058p 0 180.242p 0 180.243p 10000.0u 180.244p 0 194.306p 0 194.307p 10000.0u 194.308p 0 200.138p 0 200.139p 10000.0u 200.14p 0 202.172p 0 202.173p 10000.0u 202.174p 0 203.672p 0 203.673p 10000.0u 203.674p 0 204.638p 0 204.639p 10000.0u 204.64p 0 213.02p 0 213.021p 10000.0u 213.022p 0 223.571p 0 223.572p 10000.0u 223.573p 0 223.757p 0 223.758p 10000.0u 223.759p 0 229.211p 0 229.212p 10000.0u 229.213p 0 235.169p 0 235.17p 10000.0u 235.171p 0 253.277p 0 253.278p 10000.0u 253.279p 0 269.723p 0 269.724p 10000.0u 269.725p 0 269.756p 0 269.757p 10000.0u 269.758p 0 275.816p 0 275.817p 10000.0u 275.818p 0 280.505p 0 280.506p 10000.0u 280.507p 0 280.871p 0 280.872p 10000.0u 280.873p 0 325.04p 0 325.041p 10000.0u 325.042p 0 342.593p 0 342.594p 10000.0u 342.595p 0 343.22p 0 343.221p 10000.0u 343.222p 0 344.123p 0 344.124p 10000.0u 344.125p 0 345.971p 0 345.972p 10000.0u 345.973p 0 358.13p 0 358.131p 10000.0u 358.132p 0 362.888p 0 362.889p 10000.0u 362.89p 0 370.415p 0 370.416p 10000.0u 370.417p 0 376.469p 0 376.47p 10000.0u 376.471p 0 381.17p 0 381.171p 10000.0u 381.172p 0 396.305p 0 396.306p 10000.0u 396.307p 0 406.19p 0 406.191p 10000.0u 406.192p 0 417.341p 0 417.342p 10000.0u 417.343p 0 418.943p 0 418.944p 10000.0u 418.945p 0 431.804p 0 431.805p 10000.0u 431.806p 0 487.151p 0 487.152p 10000.0u 487.153p 0 500.687p 0 500.688p 10000.0u 500.689p 0 501.053p 0 501.054p 10000.0u 501.055p 0 523.628p 0 523.629p 10000.0u 523.63p 0 536.774p 0 536.775p 10000.0u 536.776p 0 546.689p 0 546.69p 10000.0u 546.691p 0 557.777p 0 557.778p 10000.0u 557.779p 0 569.783p 0 569.784p 10000.0u 569.785p 0 571.754p 0 571.755p 10000.0u 571.756p 0 576.704p 0 576.705p 10000.0u 576.706p 0 611.291p 0 611.292p 10000.0u 611.293p 0 615.323p 0 615.324p 10000.0u 615.325p 0 615.71p 0 615.711p 10000.0u 615.712p 0 622.004p 0 622.005p 10000.0u 622.006p 0 624.479p 0 624.48p 10000.0u 624.481p 0 665.732p 0 665.733p 10000.0u 665.734p 0 686.279p 0 686.28p 10000.0u 686.281p 0 697.526p 0 697.527p 10000.0u 697.528p 0 702.713p 0 702.714p 10000.0u 702.715p 0 704.597p 0 704.598p 10000.0u 704.599p 0 706.49p 0 706.491p 10000.0u 706.492p 0 738.908p 0 738.909p 10000.0u 738.91p 0 739.994p 0 739.995p 10000.0u 739.996p 0 764.534p 0 764.535p 10000.0u 764.536p 0 781.694p 0 781.695p 10000.0u 781.696p 0 801.278p 0 801.279p 10000.0u 801.28p 0 814.928p 0 814.929p 10000.0u 814.93p 0 822.044p 0 822.045p 10000.0u 822.046p 0 831.923p 0 831.924p 10000.0u 831.925p 0 842.492p 0 842.493p 10000.0u 842.494p 0 871.487p 0 871.488p 10000.0u 871.489p 0 872.594p 0 872.595p 10000.0u 872.596p 0 890.702p 0 890.703p 10000.0u 890.704p 0 915.434p 0 915.435p 10000.0u 915.436p 0 924.641p 0 924.642p 10000.0u 924.643p 0 927.488p 0 927.489p 10000.0u 927.49p 0 937.724p 0 937.725p 10000.0u 937.726p 0 954.599p 0 954.6p 10000.0u 954.601p 0 954.74p 0 954.741p 10000.0u 954.742p 0 969.347p 0 969.348p 10000.0u 969.349p 0 990.746p 0 990.747p 10000.0u 990.748p 0 992.324p 0 992.325p 10000.0u 992.326p 0)
IIN6 0 7 pwl(0 0 33.701p 0 33.702p 10000.0u 33.703p 0 36.263p 0 36.264p 10000.0u 36.265p 0 41.345p 0 41.346p 10000.0u 41.347p 0 49.421p 0 49.422p 10000.0u 49.423p 0 54.659p 0 54.66p 10000.0u 54.661p 0 55.796p 0 55.797p 10000.0u 55.798p 0 56.66p 0 56.661p 10000.0u 56.662p 0 73.853p 0 73.854p 10000.0u 73.855p 0 86.9p 0 86.901p 10000.0u 86.902p 0 101.342p 0 101.343p 10000.0u 101.344p 0 103.862p 0 103.863p 10000.0u 103.864p 0 115.343p 0 115.344p 10000.0u 115.345p 0 145.13p 0 145.131p 10000.0u 145.132p 0 162.287p 0 162.288p 10000.0u 162.289p 0 167.573p 0 167.574p 10000.0u 167.575p 0 167.621p 0 167.622p 10000.0u 167.623p 0 168.842p 0 168.843p 10000.0u 168.844p 0 170.888p 0 170.889p 10000.0u 170.89p 0 173.021p 0 173.022p 10000.0u 173.023p 0 180.953p 0 180.954p 10000.0u 180.955p 0 181.262p 0 181.263p 10000.0u 181.264p 0 190.586p 0 190.587p 10000.0u 190.588p 0 226.478p 0 226.479p 10000.0u 226.48p 0 229.811p 0 229.812p 10000.0u 229.813p 0 232.742p 0 232.743p 10000.0u 232.744p 0 235.205p 0 235.206p 10000.0u 235.207p 0 244.763p 0 244.764p 10000.0u 244.765p 0 274.208p 0 274.209p 10000.0u 274.21p 0 274.493p 0 274.494p 10000.0u 274.495p 0 282.857p 0 282.858p 10000.0u 282.859p 0 287.321p 0 287.322p 10000.0u 287.323p 0 322.793p 0 322.794p 10000.0u 322.795p 0 336.323p 0 336.324p 10000.0u 336.325p 0 345.053p 0 345.054p 10000.0u 345.055p 0 376.448p 0 376.449p 10000.0u 376.45p 0 377.093p 0 377.094p 10000.0u 377.095p 0 385.049p 0 385.05p 10000.0u 385.051p 0 385.991p 0 385.992p 10000.0u 385.993p 0 397.208p 0 397.209p 10000.0u 397.21p 0 397.277p 0 397.278p 10000.0u 397.279p 0 409.577p 0 409.578p 10000.0u 409.579p 0 425.765p 0 425.766p 10000.0u 425.767p 0 451.385p 0 451.386p 10000.0u 451.387p 0 455.234p 0 455.235p 10000.0u 455.236p 0 484.157p 0 484.158p 10000.0u 484.159p 0 497.942p 0 497.943p 10000.0u 497.944p 0 505.928p 0 505.929p 10000.0u 505.93p 0 511.556p 0 511.557p 10000.0u 511.558p 0 517.307p 0 517.308p 10000.0u 517.309p 0 518.228p 0 518.229p 10000.0u 518.23p 0 526.427p 0 526.428p 10000.0u 526.429p 0 529.286p 0 529.287p 10000.0u 529.288p 0 530.036p 0 530.037p 10000.0u 530.038p 0 531.704p 0 531.705p 10000.0u 531.706p 0 543.332p 0 543.333p 10000.0u 543.334p 0 551.357p 0 551.358p 10000.0u 551.359p 0 572.324p 0 572.325p 10000.0u 572.326p 0 584.441p 0 584.442p 10000.0u 584.443p 0 584.801p 0 584.802p 10000.0u 584.803p 0 589.586p 0 589.587p 10000.0u 589.588p 0 610.637p 0 610.638p 10000.0u 610.639p 0 612.008p 0 612.009p 10000.0u 612.01p 0 619.601p 0 619.602p 10000.0u 619.603p 0 633.458p 0 633.459p 10000.0u 633.46p 0 640.85p 0 640.851p 10000.0u 640.852p 0 652.889p 0 652.89p 10000.0u 652.891p 0 655.211p 0 655.212p 10000.0u 655.213p 0 657.53p 0 657.531p 10000.0u 657.532p 0 659.471p 0 659.472p 10000.0u 659.473p 0 661.496p 0 661.497p 10000.0u 661.498p 0 666.119p 0 666.12p 10000.0u 666.121p 0 676.808p 0 676.809p 10000.0u 676.81p 0 713.681p 0 713.682p 10000.0u 713.683p 0 720.146p 0 720.147p 10000.0u 720.148p 0 721.043p 0 721.044p 10000.0u 721.045p 0 730.94p 0 730.941p 10000.0u 730.942p 0 733.817p 0 733.818p 10000.0u 733.819p 0 774.209p 0 774.21p 10000.0u 774.211p 0 781.568p 0 781.569p 10000.0u 781.57p 0 783.626p 0 783.627p 10000.0u 783.628p 0 795.983p 0 795.984p 10000.0u 795.985p 0 817.634p 0 817.635p 10000.0u 817.636p 0 818.36p 0 818.361p 10000.0u 818.362p 0 821.936p 0 821.937p 10000.0u 821.938p 0 835.517p 0 835.518p 10000.0u 835.519p 0 840.431p 0 840.432p 10000.0u 840.433p 0 851.177p 0 851.178p 10000.0u 851.179p 0 860.252p 0 860.253p 10000.0u 860.254p 0 860.573p 0 860.574p 10000.0u 860.575p 0 863.957p 0 863.958p 10000.0u 863.959p 0 887.306p 0 887.307p 10000.0u 887.308p 0 920.483p 0 920.484p 10000.0u 920.485p 0 924.455p 0 924.456p 10000.0u 924.457p 0 954.209p 0 954.21p 10000.0u 954.211p 0 955.613p 0 955.614p 10000.0u 955.615p 0 968.906p 0 968.907p 10000.0u 968.908p 0 979.382p 0 979.383p 10000.0u 979.384p 0 985.193p 0 985.194p 10000.0u 985.195p 0 985.607p 0 985.608p 10000.0u 985.609p 0 986.927p 0 986.928p 10000.0u 986.929p 0 993.809p 0 993.81p 10000.0u 993.811p 0 997.931p 0 997.932p 10000.0u 997.933p 0)
IIN7 0 8 pwl(0 0 18.527p 0 18.528p 10000.0u 18.529p 0 27.578p 0 27.579p 10000.0u 27.58p 0 32.657p 0 32.658p 10000.0u 32.659p 0 33.158p 0 33.159p 10000.0u 33.16p 0 37.847p 0 37.848p 10000.0u 37.849p 0 59.855p 0 59.856p 10000.0u 59.857p 0 60.566p 0 60.567p 10000.0u 60.568p 0 68.039p 0 68.04p 10000.0u 68.041p 0 111.944p 0 111.945p 10000.0u 111.946p 0 113.444p 0 113.445p 10000.0u 113.446p 0 120.197p 0 120.198p 10000.0u 120.199p 0 136.511p 0 136.512p 10000.0u 136.513p 0 147.317p 0 147.318p 10000.0u 147.319p 0 159.068p 0 159.069p 10000.0u 159.07p 0 169.772p 0 169.773p 10000.0u 169.774p 0 176.756p 0 176.757p 10000.0u 176.758p 0 186.917p 0 186.918p 10000.0u 186.919p 0 193.631p 0 193.632p 10000.0u 193.633p 0 213.146p 0 213.147p 10000.0u 213.148p 0 216.281p 0 216.282p 10000.0u 216.283p 0 230.123p 0 230.124p 10000.0u 230.125p 0 255.458p 0 255.459p 10000.0u 255.46p 0 267.287p 0 267.288p 10000.0u 267.289p 0 276.35p 0 276.351p 10000.0u 276.352p 0 282.893p 0 282.894p 10000.0u 282.895p 0 318.311p 0 318.312p 10000.0u 318.313p 0 324.593p 0 324.594p 10000.0u 324.595p 0 324.614p 0 324.615p 10000.0u 324.616p 0 339.149p 0 339.15p 10000.0u 339.151p 0 372.236p 0 372.237p 10000.0u 372.238p 0 375.848p 0 375.849p 10000.0u 375.85p 0 375.908p 0 375.909p 10000.0u 375.91p 0 378.488p 0 378.489p 10000.0u 378.49p 0 386.579p 0 386.58p 10000.0u 386.581p 0 389.558p 0 389.559p 10000.0u 389.56p 0 399.389p 0 399.39p 10000.0u 399.391p 0 400.85p 0 400.851p 10000.0u 400.852p 0 401.168p 0 401.169p 10000.0u 401.17p 0 411.677p 0 411.678p 10000.0u 411.679p 0 428.684p 0 428.685p 10000.0u 428.686p 0 430.193p 0 430.194p 10000.0u 430.195p 0 445.985p 0 445.986p 10000.0u 445.987p 0 447.239p 0 447.24p 10000.0u 447.241p 0 458.552p 0 458.553p 10000.0u 458.554p 0 462.614p 0 462.615p 10000.0u 462.616p 0 530.18p 0 530.181p 10000.0u 530.182p 0 531.02p 0 531.021p 10000.0u 531.022p 0 534.464p 0 534.465p 10000.0u 534.466p 0 541.13p 0 541.131p 10000.0u 541.132p 0 544.748p 0 544.749p 10000.0u 544.75p 0 552.5p 0 552.501p 10000.0u 552.502p 0 554.621p 0 554.622p 10000.0u 554.623p 0 558.419p 0 558.42p 10000.0u 558.421p 0 561.959p 0 561.96p 10000.0u 561.961p 0 562.268p 0 562.269p 10000.0u 562.27p 0 573.326p 0 573.327p 10000.0u 573.328p 0 584.093p 0 584.094p 10000.0u 584.095p 0 588.257p 0 588.258p 10000.0u 588.259p 0 598.28p 0 598.281p 10000.0u 598.282p 0 603.377p 0 603.378p 10000.0u 603.379p 0 635.912p 0 635.913p 10000.0u 635.914p 0 650.963p 0 650.964p 10000.0u 650.965p 0 657.557p 0 657.558p 10000.0u 657.559p 0 675.149p 0 675.15p 10000.0u 675.151p 0 688.868p 0 688.869p 10000.0u 688.87p 0 689.501p 0 689.502p 10000.0u 689.503p 0 692.861p 0 692.862p 10000.0u 692.863p 0 702.278p 0 702.279p 10000.0u 702.28p 0 709.475p 0 709.476p 10000.0u 709.477p 0 710.888p 0 710.889p 10000.0u 710.89p 0 723.335p 0 723.336p 10000.0u 723.337p 0 728.819p 0 728.82p 10000.0u 728.821p 0 744.563p 0 744.564p 10000.0u 744.565p 0 750.83p 0 750.831p 10000.0u 750.832p 0 753.764p 0 753.765p 10000.0u 753.766p 0 759.227p 0 759.228p 10000.0u 759.229p 0 769.295p 0 769.296p 10000.0u 769.297p 0 785.411p 0 785.412p 10000.0u 785.413p 0 798.11p 0 798.111p 10000.0u 798.112p 0 801.017p 0 801.018p 10000.0u 801.019p 0 805.01p 0 805.011p 10000.0u 805.012p 0 833.153p 0 833.154p 10000.0u 833.155p 0 843.917p 0 843.918p 10000.0u 843.919p 0 846.173p 0 846.174p 10000.0u 846.175p 0 855.143p 0 855.144p 10000.0u 855.145p 0 862.667p 0 862.668p 10000.0u 862.669p 0 876.419p 0 876.42p 10000.0u 876.421p 0 886.298p 0 886.299p 10000.0u 886.3p 0 895.415p 0 895.416p 10000.0u 895.417p 0 905.573p 0 905.574p 10000.0u 905.575p 0 906.872p 0 906.873p 10000.0u 906.874p 0 907.937p 0 907.938p 10000.0u 907.939p 0 923.846p 0 923.847p 10000.0u 923.848p 0 933.806p 0 933.807p 10000.0u 933.808p 0 937.409p 0 937.41p 10000.0u 937.411p 0 939.5p 0 939.501p 10000.0u 939.502p 0 942.542p 0 942.543p 10000.0u 942.544p 0 951.32p 0 951.321p 10000.0u 951.322p 0 959.756p 0 959.757p 10000.0u 959.758p 0 961.682p 0 961.683p 10000.0u 961.684p 0 965.765p 0 965.766p 10000.0u 965.767p 0 974.615p 0 974.616p 10000.0u 974.617p 0 975.266p 0 975.267p 10000.0u 975.268p 0 975.524p 0 975.525p 10000.0u 975.526p 0 976.232p 0 976.233p 10000.0u 976.234p 0 984.146p 0 984.147p 10000.0u 984.148p 0)
IIN8 0 9 pwl(0 0 0.515p 0 0.516p 10000.0u 0.517p 0 7.115p 0 7.116p 10000.0u 7.117p 0 20.915p 0 20.916p 10000.0u 20.917p 0 21.635p 0 21.636p 10000.0u 21.637p 0 25.7p 0 25.701p 10000.0u 25.702p 0 30.794p 0 30.795p 10000.0u 30.796p 0 34.832p 0 34.833p 10000.0u 34.834p 0 50.108p 0 50.109p 10000.0u 50.11p 0 54.896p 0 54.897p 10000.0u 54.898p 0 65.84p 0 65.841p 10000.0u 65.842p 0 82.853p 0 82.854p 10000.0u 82.855p 0 87.035p 0 87.036p 10000.0u 87.037p 0 92.417p 0 92.418p 10000.0u 92.419p 0 129.779p 0 129.78p 10000.0u 129.781p 0 143.207p 0 143.208p 10000.0u 143.209p 0 144.962p 0 144.963p 10000.0u 144.964p 0 159.938p 0 159.939p 10000.0u 159.94p 0 163.217p 0 163.218p 10000.0u 163.219p 0 163.256p 0 163.257p 10000.0u 163.258p 0 166.391p 0 166.392p 10000.0u 166.393p 0 170.18p 0 170.181p 10000.0u 170.182p 0 172.511p 0 172.512p 10000.0u 172.513p 0 184.004p 0 184.005p 10000.0u 184.006p 0 212.102p 0 212.103p 10000.0u 212.104p 0 233.501p 0 233.502p 10000.0u 233.503p 0 241.634p 0 241.635p 10000.0u 241.636p 0 248.597p 0 248.598p 10000.0u 248.599p 0 254.873p 0 254.874p 10000.0u 254.875p 0 256.16p 0 256.161p 10000.0u 256.162p 0 264.422p 0 264.423p 10000.0u 264.424p 0 270.437p 0 270.438p 10000.0u 270.439p 0 272.588p 0 272.589p 10000.0u 272.59p 0 302.72p 0 302.721p 10000.0u 302.722p 0 303.149p 0 303.15p 10000.0u 303.151p 0 322.505p 0 322.506p 10000.0u 322.507p 0 329.459p 0 329.46p 10000.0u 329.461p 0 360.32p 0 360.321p 10000.0u 360.322p 0 362.471p 0 362.472p 10000.0u 362.473p 0 390.422p 0 390.423p 10000.0u 390.424p 0 400.898p 0 400.899p 10000.0u 400.9p 0 423.017p 0 423.018p 10000.0u 423.019p 0 425.879p 0 425.88p 10000.0u 425.881p 0 428.537p 0 428.538p 10000.0u 428.539p 0 443.339p 0 443.34p 10000.0u 443.341p 0 443.609p 0 443.61p 10000.0u 443.611p 0 451.535p 0 451.536p 10000.0u 451.537p 0 454.736p 0 454.737p 10000.0u 454.738p 0 461.198p 0 461.199p 10000.0u 461.2p 0 474.17p 0 474.171p 10000.0u 474.172p 0 480.461p 0 480.462p 10000.0u 480.463p 0 481.22p 0 481.221p 10000.0u 481.222p 0 483.395p 0 483.396p 10000.0u 483.397p 0 520.382p 0 520.383p 10000.0u 520.384p 0 542.807p 0 542.808p 10000.0u 542.809p 0 546.002p 0 546.003p 10000.0u 546.004p 0 557.0p 0 557.001p 10000.0u 557.002p 0 560.702p 0 560.703p 10000.0u 560.704p 0 578.939p 0 578.94p 10000.0u 578.941p 0 584.66p 0 584.661p 10000.0u 584.662p 0 589.757p 0 589.758p 10000.0u 589.759p 0 594.914p 0 594.915p 10000.0u 594.916p 0 594.947p 0 594.948p 10000.0u 594.949p 0 600.914p 0 600.915p 10000.0u 600.916p 0 604.232p 0 604.233p 10000.0u 604.234p 0 611.411p 0 611.412p 10000.0u 611.413p 0 620.864p 0 620.865p 10000.0u 620.866p 0 621.59p 0 621.591p 10000.0u 621.592p 0 635.27p 0 635.271p 10000.0u 635.272p 0 637.052p 0 637.053p 10000.0u 637.054p 0 655.982p 0 655.983p 10000.0u 655.984p 0 673.655p 0 673.656p 10000.0u 673.657p 0 688.835p 0 688.836p 10000.0u 688.837p 0 730.175p 0 730.176p 10000.0u 730.177p 0 734.435p 0 734.436p 10000.0u 734.437p 0 739.715p 0 739.716p 10000.0u 739.717p 0 742.055p 0 742.056p 10000.0u 742.057p 0 744.05p 0 744.051p 10000.0u 744.052p 0 751.34p 0 751.341p 10000.0u 751.342p 0 762.185p 0 762.186p 10000.0u 762.187p 0 800.345p 0 800.346p 10000.0u 800.347p 0 822.524p 0 822.525p 10000.0u 822.526p 0 824.747p 0 824.748p 10000.0u 824.749p 0 849.011p 0 849.012p 10000.0u 849.013p 0 855.227p 0 855.228p 10000.0u 855.229p 0 866.678p 0 866.679p 10000.0u 866.68p 0 880.328p 0 880.329p 10000.0u 880.33p 0 883.121p 0 883.122p 10000.0u 883.123p 0 894.266p 0 894.267p 10000.0u 894.268p 0 894.497p 0 894.498p 10000.0u 894.499p 0 923.303p 0 923.304p 10000.0u 923.305p 0 924.605p 0 924.606p 10000.0u 924.607p 0 929.921p 0 929.922p 10000.0u 929.923p 0 941.807p 0 941.808p 10000.0u 941.809p 0 942.263p 0 942.264p 10000.0u 942.265p 0 944.087p 0 944.088p 10000.0u 944.089p 0 952.76p 0 952.761p 10000.0u 952.762p 0 954.647p 0 954.648p 10000.0u 954.649p 0 982.241p 0 982.242p 10000.0u 982.243p 0 987.605p 0 987.606p 10000.0u 987.607p 0)
IIN9 0 10 pwl(0 0 6.959p 0 6.96p 10000.0u 6.961p 0 23.792p 0 23.793p 10000.0u 23.794p 0 33.119p 0 33.12p 10000.0u 33.121p 0 34.547p 0 34.548p 10000.0u 34.549p 0 45.071p 0 45.072p 10000.0u 45.073p 0 53.237p 0 53.238p 10000.0u 53.239p 0 53.903p 0 53.904p 10000.0u 53.905p 0 71.297p 0 71.298p 10000.0u 71.299p 0 75.935p 0 75.936p 10000.0u 75.937p 0 100.442p 0 100.443p 10000.0u 100.444p 0 112.136p 0 112.137p 10000.0u 112.138p 0 119.033p 0 119.034p 10000.0u 119.035p 0 148.256p 0 148.257p 10000.0u 148.258p 0 167.198p 0 167.199p 10000.0u 167.2p 0 167.966p 0 167.967p 10000.0u 167.968p 0 175.61p 0 175.611p 10000.0u 175.612p 0 226.121p 0 226.122p 10000.0u 226.123p 0 241.235p 0 241.236p 10000.0u 241.237p 0 248.654p 0 248.655p 10000.0u 248.656p 0 255.257p 0 255.258p 10000.0u 255.259p 0 263.462p 0 263.463p 10000.0u 263.464p 0 298.586p 0 298.587p 10000.0u 298.588p 0 348.395p 0 348.396p 10000.0u 348.397p 0 351.95p 0 351.951p 10000.0u 351.952p 0 353.96p 0 353.961p 10000.0u 353.962p 0 368.048p 0 368.049p 10000.0u 368.05p 0 395.54p 0 395.541p 10000.0u 395.542p 0 396.224p 0 396.225p 10000.0u 396.226p 0 419.54p 0 419.541p 10000.0u 419.542p 0 431.405p 0 431.406p 10000.0u 431.407p 0 436.073p 0 436.074p 10000.0u 436.075p 0 439.445p 0 439.446p 10000.0u 439.447p 0 483.857p 0 483.858p 10000.0u 483.859p 0 495.794p 0 495.795p 10000.0u 495.796p 0 501.05p 0 501.051p 10000.0u 501.052p 0 504.521p 0 504.522p 10000.0u 504.523p 0 518.471p 0 518.472p 10000.0u 518.473p 0 526.313p 0 526.314p 10000.0u 526.315p 0 529.628p 0 529.629p 10000.0u 529.63p 0 532.304p 0 532.305p 10000.0u 532.306p 0 558.716p 0 558.717p 10000.0u 558.718p 0 560.312p 0 560.313p 10000.0u 560.314p 0 562.799p 0 562.8p 10000.0u 562.801p 0 562.868p 0 562.869p 10000.0u 562.87p 0 571.571p 0 571.572p 10000.0u 571.573p 0 577.808p 0 577.809p 10000.0u 577.81p 0 579.773p 0 579.774p 10000.0u 579.775p 0 579.965p 0 579.966p 10000.0u 579.967p 0 583.721p 0 583.722p 10000.0u 583.723p 0 587.045p 0 587.046p 10000.0u 587.047p 0 590.135p 0 590.136p 10000.0u 590.137p 0 605.639p 0 605.64p 10000.0u 605.641p 0 617.258p 0 617.259p 10000.0u 617.26p 0 619.535p 0 619.536p 10000.0u 619.537p 0 629.237p 0 629.238p 10000.0u 629.239p 0 638.513p 0 638.514p 10000.0u 638.515p 0 668.492p 0 668.493p 10000.0u 668.494p 0 679.58p 0 679.581p 10000.0u 679.582p 0 694.688p 0 694.689p 10000.0u 694.69p 0 695.6p 0 695.601p 10000.0u 695.602p 0 718.751p 0 718.752p 10000.0u 718.753p 0 720.647p 0 720.648p 10000.0u 720.649p 0 736.715p 0 736.716p 10000.0u 736.717p 0 738.434p 0 738.435p 10000.0u 738.436p 0 740.528p 0 740.529p 10000.0u 740.53p 0 744.44p 0 744.441p 10000.0u 744.442p 0 754.058p 0 754.059p 10000.0u 754.06p 0 765.998p 0 765.999p 10000.0u 766.0p 0 795.923p 0 795.924p 10000.0u 795.925p 0 802.253p 0 802.254p 10000.0u 802.255p 0 814.304p 0 814.305p 10000.0u 814.306p 0 818.51p 0 818.511p 10000.0u 818.512p 0 821.27p 0 821.271p 10000.0u 821.272p 0 831.197p 0 831.198p 10000.0u 831.199p 0 864.053p 0 864.054p 10000.0u 864.055p 0 866.303p 0 866.304p 10000.0u 866.305p 0 882.467p 0 882.468p 10000.0u 882.469p 0 900.443p 0 900.444p 10000.0u 900.445p 0 921.935p 0 921.936p 10000.0u 921.937p 0 942.677p 0 942.678p 10000.0u 942.679p 0 959.963p 0 959.964p 10000.0u 959.965p 0 963.554p 0 963.555p 10000.0u 963.556p 0 979.766p 0 979.767p 10000.0u 979.768p 0 983.84p 0 983.841p 10000.0u 983.842p 0 996.194p 0 996.195p 10000.0u 996.196p 0)
IIN10 0 11 pwl(0 0 2.714p 0 2.715p 10000.0u 2.716p 0 12.218p 0 12.219p 10000.0u 12.22p 0 12.911p 0 12.912p 10000.0u 12.913p 0 44.369p 0 44.37p 10000.0u 44.371p 0 45.932p 0 45.933p 10000.0u 45.934p 0 66.101p 0 66.102p 10000.0u 66.103p 0 67.484p 0 67.485p 10000.0u 67.486p 0 71.177p 0 71.178p 10000.0u 71.179p 0 78.986p 0 78.987p 10000.0u 78.988p 0 93.488p 0 93.489p 10000.0u 93.49p 0 99.452p 0 99.453p 10000.0u 99.454p 0 113.072p 0 113.073p 10000.0u 113.074p 0 118.205p 0 118.206p 10000.0u 118.207p 0 126.719p 0 126.72p 10000.0u 126.721p 0 127.22p 0 127.221p 10000.0u 127.222p 0 138.32p 0 138.321p 10000.0u 138.322p 0 145.649p 0 145.65p 10000.0u 145.651p 0 146.348p 0 146.349p 10000.0u 146.35p 0 148.877p 0 148.878p 10000.0u 148.879p 0 171.2p 0 171.201p 10000.0u 171.202p 0 197.762p 0 197.763p 10000.0u 197.764p 0 203.258p 0 203.259p 10000.0u 203.26p 0 227.816p 0 227.817p 10000.0u 227.818p 0 236.543p 0 236.544p 10000.0u 236.545p 0 238.226p 0 238.227p 10000.0u 238.228p 0 242.177p 0 242.178p 10000.0u 242.179p 0 245.375p 0 245.376p 10000.0u 245.377p 0 258.278p 0 258.279p 10000.0u 258.28p 0 277.355p 0 277.356p 10000.0u 277.357p 0 312.122p 0 312.123p 10000.0u 312.124p 0 314.642p 0 314.643p 10000.0u 314.644p 0 315.437p 0 315.438p 10000.0u 315.439p 0 331.385p 0 331.386p 10000.0u 331.387p 0 342.182p 0 342.183p 10000.0u 342.184p 0 358.037p 0 358.038p 10000.0u 358.039p 0 365.165p 0 365.166p 10000.0u 365.167p 0 369.818p 0 369.819p 10000.0u 369.82p 0 379.253p 0 379.254p 10000.0u 379.255p 0 387.788p 0 387.789p 10000.0u 387.79p 0 392.258p 0 392.259p 10000.0u 392.26p 0 394.862p 0 394.863p 10000.0u 394.864p 0 396.056p 0 396.057p 10000.0u 396.058p 0 407.111p 0 407.112p 10000.0u 407.113p 0 416.141p 0 416.142p 10000.0u 416.143p 0 436.382p 0 436.383p 10000.0u 436.384p 0 452.18p 0 452.181p 10000.0u 452.182p 0 455.309p 0 455.31p 10000.0u 455.311p 0 469.49p 0 469.491p 10000.0u 469.492p 0 482.816p 0 482.817p 10000.0u 482.818p 0 485.6p 0 485.601p 10000.0u 485.602p 0 488.3p 0 488.301p 10000.0u 488.302p 0 499.361p 0 499.362p 10000.0u 499.363p 0 503.702p 0 503.703p 10000.0u 503.704p 0 515.762p 0 515.763p 10000.0u 515.764p 0 532.058p 0 532.059p 10000.0u 532.06p 0 541.958p 0 541.959p 10000.0u 541.96p 0 551.987p 0 551.988p 10000.0u 551.989p 0 559.28p 0 559.281p 10000.0u 559.282p 0 563.573p 0 563.574p 10000.0u 563.575p 0 564.233p 0 564.234p 10000.0u 564.235p 0 569.198p 0 569.199p 10000.0u 569.2p 0 584.999p 0 585.0p 10000.0u 585.001p 0 590.882p 0 590.883p 10000.0u 590.884p 0 592.811p 0 592.812p 10000.0u 592.813p 0 603.242p 0 603.243p 10000.0u 603.244p 0 614.567p 0 614.568p 10000.0u 614.569p 0 617.414p 0 617.415p 10000.0u 617.416p 0 628.256p 0 628.257p 10000.0u 628.258p 0 631.934p 0 631.935p 10000.0u 631.936p 0 645.458p 0 645.459p 10000.0u 645.46p 0 664.175p 0 664.176p 10000.0u 664.177p 0 664.952p 0 664.953p 10000.0u 664.954p 0 666.575p 0 666.576p 10000.0u 666.577p 0 684.26p 0 684.261p 10000.0u 684.262p 0 686.663p 0 686.664p 10000.0u 686.665p 0 691.328p 0 691.329p 10000.0u 691.33p 0 693.92p 0 693.921p 10000.0u 693.922p 0 703.628p 0 703.629p 10000.0u 703.63p 0 703.715p 0 703.716p 10000.0u 703.717p 0 713.78p 0 713.781p 10000.0u 713.782p 0 722.687p 0 722.688p 10000.0u 722.689p 0 756.749p 0 756.75p 10000.0u 756.751p 0 757.739p 0 757.74p 10000.0u 757.741p 0 761.087p 0 761.088p 10000.0u 761.089p 0 761.192p 0 761.193p 10000.0u 761.194p 0 762.05p 0 762.051p 10000.0u 762.052p 0 777.686p 0 777.687p 10000.0u 777.688p 0 796.607p 0 796.608p 10000.0u 796.609p 0 800.792p 0 800.793p 10000.0u 800.794p 0 810.464p 0 810.465p 10000.0u 810.466p 0 815.018p 0 815.019p 10000.0u 815.02p 0 834.605p 0 834.606p 10000.0u 834.607p 0 855.38p 0 855.381p 10000.0u 855.382p 0 860.978p 0 860.979p 10000.0u 860.98p 0 861.095p 0 861.096p 10000.0u 861.097p 0 868.871p 0 868.872p 10000.0u 868.873p 0 874.934p 0 874.935p 10000.0u 874.936p 0 875.393p 0 875.394p 10000.0u 875.395p 0 876.797p 0 876.798p 10000.0u 876.799p 0 878.99p 0 878.991p 10000.0u 878.992p 0 888.998p 0 888.999p 10000.0u 889.0p 0 898.607p 0 898.608p 10000.0u 898.609p 0 900.572p 0 900.573p 10000.0u 900.574p 0 902.213p 0 902.214p 10000.0u 902.215p 0 951.134p 0 951.135p 10000.0u 951.136p 0 955.151p 0 955.152p 10000.0u 955.153p 0 965.123p 0 965.124p 10000.0u 965.125p 0 966.182p 0 966.183p 10000.0u 966.184p 0 968.135p 0 968.136p 10000.0u 968.137p 0 968.273p 0 968.274p 10000.0u 968.275p 0 972.455p 0 972.456p 10000.0u 972.457p 0 982.886p 0 982.887p 10000.0u 982.888p 0 990.152p 0 990.153p 10000.0u 990.154p 0)
IIN11 0 12 pwl(0 0 3.863p 0 3.864p 10000.0u 3.865p 0 12.254p 0 12.255p 10000.0u 12.256p 0 29.24p 0 29.241p 10000.0u 29.242p 0 74.498p 0 74.499p 10000.0u 74.5p 0 99.692p 0 99.693p 10000.0u 99.694p 0 114.761p 0 114.762p 10000.0u 114.763p 0 115.409p 0 115.41p 10000.0u 115.411p 0 137.237p 0 137.238p 10000.0u 137.239p 0 137.645p 0 137.646p 10000.0u 137.647p 0 138.605p 0 138.606p 10000.0u 138.607p 0 173.198p 0 173.199p 10000.0u 173.2p 0 186.527p 0 186.528p 10000.0u 186.529p 0 188.135p 0 188.136p 10000.0u 188.137p 0 189.722p 0 189.723p 10000.0u 189.724p 0 191.123p 0 191.124p 10000.0u 191.125p 0 191.927p 0 191.928p 10000.0u 191.929p 0 206.759p 0 206.76p 10000.0u 206.761p 0 219.371p 0 219.372p 10000.0u 219.373p 0 220.559p 0 220.56p 10000.0u 220.561p 0 236.39p 0 236.391p 10000.0u 236.392p 0 241.643p 0 241.644p 10000.0u 241.645p 0 243.482p 0 243.483p 10000.0u 243.484p 0 245.711p 0 245.712p 10000.0u 245.713p 0 247.7p 0 247.701p 10000.0u 247.702p 0 268.409p 0 268.41p 10000.0u 268.411p 0 283.046p 0 283.047p 10000.0u 283.048p 0 285.647p 0 285.648p 10000.0u 285.649p 0 290.981p 0 290.982p 10000.0u 290.983p 0 291.746p 0 291.747p 10000.0u 291.748p 0 301.64p 0 301.641p 10000.0u 301.642p 0 303.218p 0 303.219p 10000.0u 303.22p 0 308.987p 0 308.988p 10000.0u 308.989p 0 332.996p 0 332.997p 10000.0u 332.998p 0 353.048p 0 353.049p 10000.0u 353.05p 0 354.191p 0 354.192p 10000.0u 354.193p 0 370.523p 0 370.524p 10000.0u 370.525p 0 371.444p 0 371.445p 10000.0u 371.446p 0 380.624p 0 380.625p 10000.0u 380.626p 0 397.652p 0 397.653p 10000.0u 397.654p 0 402.818p 0 402.819p 10000.0u 402.82p 0 408.5p 0 408.501p 10000.0u 408.502p 0 413.825p 0 413.826p 10000.0u 413.827p 0 422.813p 0 422.814p 10000.0u 422.815p 0 432.848p 0 432.849p 10000.0u 432.85p 0 442.286p 0 442.287p 10000.0u 442.288p 0 456.743p 0 456.744p 10000.0u 456.745p 0 494.732p 0 494.733p 10000.0u 494.734p 0 497.846p 0 497.847p 10000.0u 497.848p 0 543.383p 0 543.384p 10000.0u 543.385p 0 549.713p 0 549.714p 10000.0u 549.715p 0 550.109p 0 550.11p 10000.0u 550.111p 0 557.291p 0 557.292p 10000.0u 557.293p 0 559.001p 0 559.002p 10000.0u 559.003p 0 559.592p 0 559.593p 10000.0u 559.594p 0 562.232p 0 562.233p 10000.0u 562.234p 0 600.206p 0 600.207p 10000.0u 600.208p 0 605.234p 0 605.235p 10000.0u 605.236p 0 606.602p 0 606.603p 10000.0u 606.604p 0 609.584p 0 609.585p 10000.0u 609.586p 0 628.649p 0 628.65p 10000.0u 628.651p 0 636.602p 0 636.603p 10000.0u 636.604p 0 644.996p 0 644.997p 10000.0u 644.998p 0 647.249p 0 647.25p 10000.0u 647.251p 0 647.39p 0 647.391p 10000.0u 647.392p 0 654.803p 0 654.804p 10000.0u 654.805p 0 657.08p 0 657.081p 10000.0u 657.082p 0 664.745p 0 664.746p 10000.0u 664.747p 0 673.715p 0 673.716p 10000.0u 673.717p 0 678.461p 0 678.462p 10000.0u 678.463p 0 709.646p 0 709.647p 10000.0u 709.648p 0 733.433p 0 733.434p 10000.0u 733.435p 0 758.393p 0 758.394p 10000.0u 758.395p 0 768.674p 0 768.675p 10000.0u 768.676p 0 771.851p 0 771.852p 10000.0u 771.853p 0 778.382p 0 778.383p 10000.0u 778.384p 0 779.003p 0 779.004p 10000.0u 779.005p 0 794.405p 0 794.406p 10000.0u 794.407p 0 819.305p 0 819.306p 10000.0u 819.307p 0 825.419p 0 825.42p 10000.0u 825.421p 0 832.457p 0 832.458p 10000.0u 832.459p 0 833.894p 0 833.895p 10000.0u 833.896p 0 840.506p 0 840.507p 10000.0u 840.508p 0 852.722p 0 852.723p 10000.0u 852.724p 0 876.809p 0 876.81p 10000.0u 876.811p 0 877.052p 0 877.053p 10000.0u 877.054p 0 882.164p 0 882.165p 10000.0u 882.166p 0 882.26p 0 882.261p 10000.0u 882.262p 0 884.186p 0 884.187p 10000.0u 884.188p 0 887.165p 0 887.166p 10000.0u 887.167p 0 890.858p 0 890.859p 10000.0u 890.86p 0 892.805p 0 892.806p 10000.0u 892.807p 0 908.27p 0 908.271p 10000.0u 908.272p 0 914.9p 0 914.901p 10000.0u 914.902p 0 926.435p 0 926.436p 10000.0u 926.437p 0 927.515p 0 927.516p 10000.0u 927.517p 0 948.857p 0 948.858p 10000.0u 948.859p 0 952.43p 0 952.431p 10000.0u 952.432p 0 954.302p 0 954.303p 10000.0u 954.304p 0 954.425p 0 954.426p 10000.0u 954.427p 0 968.648p 0 968.649p 10000.0u 968.65p 0 975.059p 0 975.06p 10000.0u 975.061p 0 984.203p 0 984.204p 10000.0u 984.205p 0 985.886p 0 985.887p 10000.0u 985.888p 0 997.979p 0 997.98p 10000.0u 997.981p 0 998.897p 0 998.898p 10000.0u 998.899p 0)
IIN12 0 13 pwl(0 0 1.97p 0 1.971p 10000.0u 1.972p 0 43.376p 0 43.377p 10000.0u 43.378p 0 43.784p 0 43.785p 10000.0u 43.786p 0 67.901p 0 67.902p 10000.0u 67.903p 0 75.941p 0 75.942p 10000.0u 75.943p 0 79.67p 0 79.671p 10000.0u 79.672p 0 94.34p 0 94.341p 10000.0u 94.342p 0 112.703p 0 112.704p 10000.0u 112.705p 0 122.789p 0 122.79p 10000.0u 122.791p 0 130.067p 0 130.068p 10000.0u 130.069p 0 138.878p 0 138.879p 10000.0u 138.88p 0 159.92p 0 159.921p 10000.0u 159.922p 0 167.51p 0 167.511p 10000.0u 167.512p 0 169.181p 0 169.182p 10000.0u 169.183p 0 219.959p 0 219.96p 10000.0u 219.961p 0 224.342p 0 224.343p 10000.0u 224.344p 0 244.235p 0 244.236p 10000.0u 244.237p 0 262.7p 0 262.701p 10000.0u 262.702p 0 282.122p 0 282.123p 10000.0u 282.124p 0 282.932p 0 282.933p 10000.0u 282.934p 0 285.278p 0 285.279p 10000.0u 285.28p 0 312.041p 0 312.042p 10000.0u 312.043p 0 359.663p 0 359.664p 10000.0u 359.665p 0 370.484p 0 370.485p 10000.0u 370.486p 0 382.172p 0 382.173p 10000.0u 382.174p 0 404.087p 0 404.088p 10000.0u 404.089p 0 409.718p 0 409.719p 10000.0u 409.72p 0 424.367p 0 424.368p 10000.0u 424.369p 0 428.945p 0 428.946p 10000.0u 428.947p 0 429.554p 0 429.555p 10000.0u 429.556p 0 433.925p 0 433.926p 10000.0u 433.927p 0 435.095p 0 435.096p 10000.0u 435.097p 0 441.23p 0 441.231p 10000.0u 441.232p 0 444.809p 0 444.81p 10000.0u 444.811p 0 445.544p 0 445.545p 10000.0u 445.546p 0 457.673p 0 457.674p 10000.0u 457.675p 0 459.5p 0 459.501p 10000.0u 459.502p 0 460.805p 0 460.806p 10000.0u 460.807p 0 470.678p 0 470.679p 10000.0u 470.68p 0 477.791p 0 477.792p 10000.0u 477.793p 0 525.128p 0 525.129p 10000.0u 525.13p 0 526.7p 0 526.701p 10000.0u 526.702p 0 536.504p 0 536.505p 10000.0u 536.506p 0 567.059p 0 567.06p 10000.0u 567.061p 0 613.748p 0 613.749p 10000.0u 613.75p 0 617.591p 0 617.592p 10000.0u 617.593p 0 654.596p 0 654.597p 10000.0u 654.598p 0 664.232p 0 664.233p 10000.0u 664.234p 0 688.598p 0 688.599p 10000.0u 688.6p 0 688.664p 0 688.665p 10000.0u 688.666p 0 691.208p 0 691.209p 10000.0u 691.21p 0 695.795p 0 695.796p 10000.0u 695.797p 0 700.16p 0 700.161p 10000.0u 700.162p 0 703.133p 0 703.134p 10000.0u 703.135p 0 705.008p 0 705.009p 10000.0u 705.01p 0 722.579p 0 722.58p 10000.0u 722.581p 0 723.341p 0 723.342p 10000.0u 723.343p 0 732.608p 0 732.609p 10000.0u 732.61p 0 734.264p 0 734.265p 10000.0u 734.266p 0 743.798p 0 743.799p 10000.0u 743.8p 0 757.7p 0 757.701p 10000.0u 757.702p 0 788.306p 0 788.307p 10000.0u 788.308p 0 820.292p 0 820.293p 10000.0u 820.294p 0 833.252p 0 833.253p 10000.0u 833.254p 0 856.826p 0 856.827p 10000.0u 856.828p 0 868.934p 0 868.935p 10000.0u 868.936p 0 872.147p 0 872.148p 10000.0u 872.149p 0 876.968p 0 876.969p 10000.0u 876.97p 0 913.883p 0 913.884p 10000.0u 913.885p 0 929.057p 0 929.058p 10000.0u 929.059p 0 976.676p 0 976.677p 10000.0u 976.678p 0 981.464p 0 981.465p 10000.0u 981.466p 0 985.016p 0 985.017p 10000.0u 985.018p 0 989.417p 0 989.418p 10000.0u 989.419p 0 990.818p 0 990.819p 10000.0u 990.82p 0)
IIN13 0 14 pwl(0 0 3.416p 0 3.417p 10000.0u 3.418p 0 15.044p 0 15.045p 10000.0u 15.046p 0 16.508p 0 16.509p 10000.0u 16.51p 0 22.121p 0 22.122p 10000.0u 22.123p 0 23.564p 0 23.565p 10000.0u 23.566p 0 29.642p 0 29.643p 10000.0u 29.644p 0 31.586p 0 31.587p 10000.0u 31.588p 0 35.195p 0 35.196p 10000.0u 35.197p 0 39.398p 0 39.399p 10000.0u 39.4p 0 39.407p 0 39.408p 10000.0u 39.409p 0 51.062p 0 51.063p 10000.0u 51.064p 0 66.482p 0 66.483p 10000.0u 66.484p 0 66.542p 0 66.543p 10000.0u 66.544p 0 70.745p 0 70.746p 10000.0u 70.747p 0 109.166p 0 109.167p 10000.0u 109.168p 0 129.308p 0 129.309p 10000.0u 129.31p 0 131.753p 0 131.754p 10000.0u 131.755p 0 133.589p 0 133.59p 10000.0u 133.591p 0 137.393p 0 137.394p 10000.0u 137.395p 0 149.036p 0 149.037p 10000.0u 149.038p 0 164.024p 0 164.025p 10000.0u 164.026p 0 174.761p 0 174.762p 10000.0u 174.763p 0 194.015p 0 194.016p 10000.0u 194.017p 0 205.931p 0 205.932p 10000.0u 205.933p 0 206.45p 0 206.451p 10000.0u 206.452p 0 206.885p 0 206.886p 10000.0u 206.887p 0 207.971p 0 207.972p 10000.0u 207.973p 0 212.507p 0 212.508p 10000.0u 212.509p 0 216.143p 0 216.144p 10000.0u 216.145p 0 219.101p 0 219.102p 10000.0u 219.103p 0 225.611p 0 225.612p 10000.0u 225.613p 0 227.252p 0 227.253p 10000.0u 227.254p 0 236.699p 0 236.7p 10000.0u 236.701p 0 243.431p 0 243.432p 10000.0u 243.433p 0 265.025p 0 265.026p 10000.0u 265.027p 0 283.52p 0 283.521p 10000.0u 283.522p 0 286.484p 0 286.485p 10000.0u 286.486p 0 303.218p 0 303.219p 10000.0u 303.22p 0 316.181p 0 316.182p 10000.0u 316.183p 0 319.034p 0 319.035p 10000.0u 319.036p 0 320.612p 0 320.613p 10000.0u 320.614p 0 322.673p 0 322.674p 10000.0u 322.675p 0 325.76p 0 325.761p 10000.0u 325.762p 0 328.829p 0 328.83p 10000.0u 328.831p 0 341.495p 0 341.496p 10000.0u 341.497p 0 352.769p 0 352.77p 10000.0u 352.771p 0 367.028p 0 367.029p 10000.0u 367.03p 0 394.712p 0 394.713p 10000.0u 394.714p 0 402.689p 0 402.69p 10000.0u 402.691p 0 402.836p 0 402.837p 10000.0u 402.838p 0 402.962p 0 402.963p 10000.0u 402.964p 0 407.864p 0 407.865p 10000.0u 407.866p 0 420.344p 0 420.345p 10000.0u 420.346p 0 443.993p 0 443.994p 10000.0u 443.995p 0 454.796p 0 454.797p 10000.0u 454.798p 0 488.363p 0 488.364p 10000.0u 488.365p 0 509.624p 0 509.625p 10000.0u 509.626p 0 511.955p 0 511.956p 10000.0u 511.957p 0 512.075p 0 512.076p 10000.0u 512.077p 0 532.328p 0 532.329p 10000.0u 532.33p 0 534.614p 0 534.615p 10000.0u 534.616p 0 535.16p 0 535.161p 10000.0u 535.162p 0 547.337p 0 547.338p 10000.0u 547.339p 0 559.664p 0 559.665p 10000.0u 559.666p 0 567.347p 0 567.348p 10000.0u 567.349p 0 569.819p 0 569.82p 10000.0u 569.821p 0 571.958p 0 571.959p 10000.0u 571.96p 0 573.413p 0 573.414p 10000.0u 573.415p 0 589.262p 0 589.263p 10000.0u 589.264p 0 609.872p 0 609.873p 10000.0u 609.874p 0 627.11p 0 627.111p 10000.0u 627.112p 0 637.085p 0 637.086p 10000.0u 637.087p 0 653.495p 0 653.496p 10000.0u 653.497p 0 660.707p 0 660.708p 10000.0u 660.709p 0 666.491p 0 666.492p 10000.0u 666.493p 0 694.343p 0 694.344p 10000.0u 694.345p 0 705.2p 0 705.201p 10000.0u 705.202p 0 707.654p 0 707.655p 10000.0u 707.656p 0 709.28p 0 709.281p 10000.0u 709.282p 0 712.499p 0 712.5p 10000.0u 712.501p 0 753.041p 0 753.042p 10000.0u 753.043p 0 758.774p 0 758.775p 10000.0u 758.776p 0 768.419p 0 768.42p 10000.0u 768.421p 0 776.924p 0 776.925p 10000.0u 776.926p 0 780.224p 0 780.225p 10000.0u 780.226p 0 828.875p 0 828.876p 10000.0u 828.877p 0 828.959p 0 828.96p 10000.0u 828.961p 0 848.339p 0 848.34p 10000.0u 848.341p 0 851.498p 0 851.499p 10000.0u 851.5p 0 871.202p 0 871.203p 10000.0u 871.204p 0 872.951p 0 872.952p 10000.0u 872.953p 0 876.677p 0 876.678p 10000.0u 876.679p 0 881.561p 0 881.562p 10000.0u 881.563p 0 881.579p 0 881.58p 10000.0u 881.581p 0 896.279p 0 896.28p 10000.0u 896.281p 0 910.505p 0 910.506p 10000.0u 910.507p 0 912.116p 0 912.117p 10000.0u 912.118p 0 920.357p 0 920.358p 10000.0u 920.359p 0 928.823p 0 928.824p 10000.0u 928.825p 0 957.392p 0 957.393p 10000.0u 957.394p 0 985.253p 0 985.254p 10000.0u 985.255p 0 995.732p 0 995.733p 10000.0u 995.734p 0 996.677p 0 996.678p 10000.0u 996.679p 0)
IIN14 0 15 pwl(0 0 0.338p 0 0.339p 10000.0u 0.34p 0 18.563p 0 18.564p 10000.0u 18.565p 0 32.672p 0 32.673p 10000.0u 32.674p 0 51.401p 0 51.402p 10000.0u 51.403p 0 57.347p 0 57.348p 10000.0u 57.349p 0 64.271p 0 64.272p 10000.0u 64.273p 0 70.019p 0 70.02p 10000.0u 70.021p 0 88.268p 0 88.269p 10000.0u 88.27p 0 100.508p 0 100.509p 10000.0u 100.51p 0 102.953p 0 102.954p 10000.0u 102.955p 0 108.119p 0 108.12p 10000.0u 108.121p 0 137.756p 0 137.757p 10000.0u 137.758p 0 146.348p 0 146.349p 10000.0u 146.35p 0 151.79p 0 151.791p 10000.0u 151.792p 0 156.548p 0 156.549p 10000.0u 156.55p 0 184.25p 0 184.251p 10000.0u 184.252p 0 188.252p 0 188.253p 10000.0u 188.254p 0 211.604p 0 211.605p 10000.0u 211.606p 0 212.582p 0 212.583p 10000.0u 212.584p 0 224.045p 0 224.046p 10000.0u 224.047p 0 226.271p 0 226.272p 10000.0u 226.273p 0 228.386p 0 228.387p 10000.0u 228.388p 0 233.969p 0 233.97p 10000.0u 233.971p 0 238.634p 0 238.635p 10000.0u 238.636p 0 241.31p 0 241.311p 10000.0u 241.312p 0 243.047p 0 243.048p 10000.0u 243.049p 0 243.41p 0 243.411p 10000.0u 243.412p 0 247.271p 0 247.272p 10000.0u 247.273p 0 269.972p 0 269.973p 10000.0u 269.974p 0 270.452p 0 270.453p 10000.0u 270.454p 0 273.173p 0 273.174p 10000.0u 273.175p 0 293.372p 0 293.373p 10000.0u 293.374p 0 299.723p 0 299.724p 10000.0u 299.725p 0 308.162p 0 308.163p 10000.0u 308.164p 0 310.325p 0 310.326p 10000.0u 310.327p 0 313.364p 0 313.365p 10000.0u 313.366p 0 314.735p 0 314.736p 10000.0u 314.737p 0 331.118p 0 331.119p 10000.0u 331.12p 0 342.842p 0 342.843p 10000.0u 342.844p 0 367.817p 0 367.818p 10000.0u 367.819p 0 370.652p 0 370.653p 10000.0u 370.654p 0 378.998p 0 378.999p 10000.0u 379.0p 0 390.869p 0 390.87p 10000.0u 390.871p 0 408.878p 0 408.879p 10000.0u 408.88p 0 416.822p 0 416.823p 10000.0u 416.824p 0 424.334p 0 424.335p 10000.0u 424.336p 0 444.926p 0 444.927p 10000.0u 444.928p 0 451.352p 0 451.353p 10000.0u 451.354p 0 453.326p 0 453.327p 10000.0u 453.328p 0 458.669p 0 458.67p 10000.0u 458.671p 0 459.239p 0 459.24p 10000.0u 459.241p 0 467.222p 0 467.223p 10000.0u 467.224p 0 468.251p 0 468.252p 10000.0u 468.253p 0 498.596p 0 498.597p 10000.0u 498.598p 0 506.747p 0 506.748p 10000.0u 506.749p 0 514.565p 0 514.566p 10000.0u 514.567p 0 516.962p 0 516.963p 10000.0u 516.964p 0 526.748p 0 526.749p 10000.0u 526.75p 0 538.094p 0 538.095p 10000.0u 538.096p 0 553.37p 0 553.371p 10000.0u 553.372p 0 554.597p 0 554.598p 10000.0u 554.599p 0 575.486p 0 575.487p 10000.0u 575.488p 0 587.006p 0 587.007p 10000.0u 587.008p 0 597.359p 0 597.36p 10000.0u 597.361p 0 607.424p 0 607.425p 10000.0u 607.426p 0 609.197p 0 609.198p 10000.0u 609.199p 0 614.51p 0 614.511p 10000.0u 614.512p 0 621.884p 0 621.885p 10000.0u 621.886p 0 657.419p 0 657.42p 10000.0u 657.421p 0 661.745p 0 661.746p 10000.0u 661.747p 0 698.567p 0 698.568p 10000.0u 698.569p 0 702.491p 0 702.492p 10000.0u 702.493p 0 707.465p 0 707.466p 10000.0u 707.467p 0 710.597p 0 710.598p 10000.0u 710.599p 0 723.014p 0 723.015p 10000.0u 723.016p 0 732.737p 0 732.738p 10000.0u 732.739p 0 754.178p 0 754.179p 10000.0u 754.18p 0 759.941p 0 759.942p 10000.0u 759.943p 0 766.154p 0 766.155p 10000.0u 766.156p 0 787.484p 0 787.485p 10000.0u 787.486p 0 794.015p 0 794.016p 10000.0u 794.017p 0 798.392p 0 798.393p 10000.0u 798.394p 0 803.006p 0 803.007p 10000.0u 803.008p 0 803.03p 0 803.031p 10000.0u 803.032p 0 827.78p 0 827.781p 10000.0u 827.782p 0 846.131p 0 846.132p 10000.0u 846.133p 0 846.821p 0 846.822p 10000.0u 846.823p 0 877.286p 0 877.287p 10000.0u 877.288p 0 878.339p 0 878.34p 10000.0u 878.341p 0 881.774p 0 881.775p 10000.0u 881.776p 0 892.826p 0 892.827p 10000.0u 892.828p 0 896.54p 0 896.541p 10000.0u 896.542p 0 901.673p 0 901.674p 10000.0u 901.675p 0 909.809p 0 909.81p 10000.0u 909.811p 0 909.941p 0 909.942p 10000.0u 909.943p 0 911.873p 0 911.874p 10000.0u 911.875p 0 924.323p 0 924.324p 10000.0u 924.325p 0 936.116p 0 936.117p 10000.0u 936.118p 0 936.869p 0 936.87p 10000.0u 936.871p 0 947.984p 0 947.985p 10000.0u 947.986p 0 958.577p 0 958.578p 10000.0u 958.579p 0 965.195p 0 965.196p 10000.0u 965.197p 0 973.004p 0 973.005p 10000.0u 973.006p 0 977.93p 0 977.931p 10000.0u 977.932p 0 978.287p 0 978.288p 10000.0u 978.289p 0 978.611p 0 978.612p 10000.0u 978.613p 0 979.637p 0 979.638p 10000.0u 979.639p 0 983.939p 0 983.94p 10000.0u 983.941p 0)
IIN15 0 16 pwl(0 0 0.731p 0 0.732p 10000.0u 0.733p 0 12.809p 0 12.81p 10000.0u 12.811p 0 15.164p 0 15.165p 10000.0u 15.166p 0 16.217p 0 16.218p 10000.0u 16.219p 0 57.293p 0 57.294p 10000.0u 57.295p 0 58.94p 0 58.941p 10000.0u 58.942p 0 67.436p 0 67.437p 10000.0u 67.438p 0 94.973p 0 94.974p 10000.0u 94.975p 0 112.625p 0 112.626p 10000.0u 112.627p 0 115.052p 0 115.053p 10000.0u 115.054p 0 130.211p 0 130.212p 10000.0u 130.213p 0 143.15p 0 143.151p 10000.0u 143.152p 0 149.753p 0 149.754p 10000.0u 149.755p 0 156.383p 0 156.384p 10000.0u 156.385p 0 157.043p 0 157.044p 10000.0u 157.045p 0 159.887p 0 159.888p 10000.0u 159.889p 0 160.268p 0 160.269p 10000.0u 160.27p 0 177.341p 0 177.342p 10000.0u 177.343p 0 179.243p 0 179.244p 10000.0u 179.245p 0 181.43p 0 181.431p 10000.0u 181.432p 0 187.289p 0 187.29p 10000.0u 187.291p 0 190.403p 0 190.404p 10000.0u 190.405p 0 191.201p 0 191.202p 10000.0u 191.203p 0 214.394p 0 214.395p 10000.0u 214.396p 0 229.538p 0 229.539p 10000.0u 229.54p 0 231.821p 0 231.822p 10000.0u 231.823p 0 252.443p 0 252.444p 10000.0u 252.445p 0 265.304p 0 265.305p 10000.0u 265.306p 0 265.91p 0 265.911p 10000.0u 265.912p 0 272.111p 0 272.112p 10000.0u 272.113p 0 293.795p 0 293.796p 10000.0u 293.797p 0 302.939p 0 302.94p 10000.0u 302.941p 0 314.777p 0 314.778p 10000.0u 314.779p 0 328.898p 0 328.899p 10000.0u 328.9p 0 352.679p 0 352.68p 10000.0u 352.681p 0 376.133p 0 376.134p 10000.0u 376.135p 0 377.423p 0 377.424p 10000.0u 377.425p 0 384.296p 0 384.297p 10000.0u 384.298p 0 396.221p 0 396.222p 10000.0u 396.223p 0 399.641p 0 399.642p 10000.0u 399.643p 0 408.749p 0 408.75p 10000.0u 408.751p 0 428.027p 0 428.028p 10000.0u 428.029p 0 442.676p 0 442.677p 10000.0u 442.678p 0 456.998p 0 456.999p 10000.0u 457.0p 0 470.879p 0 470.88p 10000.0u 470.881p 0 478.139p 0 478.14p 10000.0u 478.141p 0 493.043p 0 493.044p 10000.0u 493.045p 0 505.547p 0 505.548p 10000.0u 505.549p 0 506.429p 0 506.43p 10000.0u 506.431p 0 513.998p 0 513.999p 10000.0u 514.0p 0 526.439p 0 526.44p 10000.0u 526.441p 0 527.744p 0 527.745p 10000.0u 527.746p 0 540.767p 0 540.768p 10000.0u 540.769p 0 559.544p 0 559.545p 10000.0u 559.546p 0 559.589p 0 559.59p 10000.0u 559.591p 0 570.836p 0 570.837p 10000.0u 570.838p 0 572.045p 0 572.046p 10000.0u 572.047p 0 583.268p 0 583.269p 10000.0u 583.27p 0 606.53p 0 606.531p 10000.0u 606.532p 0 608.837p 0 608.838p 10000.0u 608.839p 0 619.82p 0 619.821p 10000.0u 619.822p 0 624.818p 0 624.819p 10000.0u 624.82p 0 625.568p 0 625.569p 10000.0u 625.57p 0 626.489p 0 626.49p 10000.0u 626.491p 0 628.115p 0 628.116p 10000.0u 628.117p 0 631.262p 0 631.263p 10000.0u 631.264p 0 632.657p 0 632.658p 10000.0u 632.659p 0 649.862p 0 649.863p 10000.0u 649.864p 0 658.589p 0 658.59p 10000.0u 658.591p 0 659.963p 0 659.964p 10000.0u 659.965p 0 674.252p 0 674.253p 10000.0u 674.254p 0 676.931p 0 676.932p 10000.0u 676.933p 0 709.454p 0 709.455p 10000.0u 709.456p 0 713.825p 0 713.826p 10000.0u 713.827p 0 720.917p 0 720.918p 10000.0u 720.919p 0 720.971p 0 720.972p 10000.0u 720.973p 0 721.517p 0 721.518p 10000.0u 721.519p 0 726.299p 0 726.3p 10000.0u 726.301p 0 730.733p 0 730.734p 10000.0u 730.735p 0 736.697p 0 736.698p 10000.0u 736.699p 0 756.131p 0 756.132p 10000.0u 756.133p 0 776.504p 0 776.505p 10000.0u 776.506p 0 779.216p 0 779.217p 10000.0u 779.218p 0 810.614p 0 810.615p 10000.0u 810.616p 0 814.304p 0 814.305p 10000.0u 814.306p 0 827.492p 0 827.493p 10000.0u 827.494p 0 840.5p 0 840.501p 10000.0u 840.502p 0 851.378p 0 851.379p 10000.0u 851.38p 0 858.812p 0 858.813p 10000.0u 858.814p 0 860.909p 0 860.91p 10000.0u 860.911p 0 871.28p 0 871.281p 10000.0u 871.282p 0 874.79p 0 874.791p 10000.0u 874.792p 0 915.293p 0 915.294p 10000.0u 915.295p 0 920.927p 0 920.928p 10000.0u 920.929p 0 945.788p 0 945.789p 10000.0u 945.79p 0 992.075p 0 992.076p 10000.0u 992.077p 0 992.135p 0 992.136p 10000.0u 992.137p 0 994.316p 0 994.317p 10000.0u 994.318p 0 996.434p 0 996.435p 10000.0u 996.436p 0)
IIN16 0 17 pwl(0 0 14.924p 0 14.925p 10000.0u 14.926p 0 21.455p 0 21.456p 10000.0u 21.457p 0 23.525p 0 23.526p 10000.0u 23.527p 0 26.18p 0 26.181p 10000.0u 26.182p 0 32.27p 0 32.271p 10000.0u 32.272p 0 35.996p 0 35.997p 10000.0u 35.998p 0 41.669p 0 41.67p 10000.0u 41.671p 0 60.752p 0 60.753p 10000.0u 60.754p 0 64.934p 0 64.935p 10000.0u 64.936p 0 77.942p 0 77.943p 10000.0u 77.944p 0 89.237p 0 89.238p 10000.0u 89.239p 0 94.445p 0 94.446p 10000.0u 94.447p 0 111.002p 0 111.003p 10000.0u 111.004p 0 115.862p 0 115.863p 10000.0u 115.864p 0 123.605p 0 123.606p 10000.0u 123.607p 0 128.555p 0 128.556p 10000.0u 128.557p 0 129.419p 0 129.42p 10000.0u 129.421p 0 136.853p 0 136.854p 10000.0u 136.855p 0 157.43p 0 157.431p 10000.0u 157.432p 0 166.646p 0 166.647p 10000.0u 166.648p 0 183.629p 0 183.63p 10000.0u 183.631p 0 186.743p 0 186.744p 10000.0u 186.745p 0 189.875p 0 189.876p 10000.0u 189.877p 0 200.375p 0 200.376p 10000.0u 200.377p 0 203.384p 0 203.385p 10000.0u 203.386p 0 204.746p 0 204.747p 10000.0u 204.748p 0 209.159p 0 209.16p 10000.0u 209.161p 0 214.148p 0 214.149p 10000.0u 214.15p 0 232.199p 0 232.2p 10000.0u 232.201p 0 275.498p 0 275.499p 10000.0u 275.5p 0 279.593p 0 279.594p 10000.0u 279.595p 0 282.908p 0 282.909p 10000.0u 282.91p 0 302.501p 0 302.502p 10000.0u 302.503p 0 312.308p 0 312.309p 10000.0u 312.31p 0 327.581p 0 327.582p 10000.0u 327.583p 0 327.914p 0 327.915p 10000.0u 327.916p 0 337.475p 0 337.476p 10000.0u 337.477p 0 339.122p 0 339.123p 10000.0u 339.124p 0 354.278p 0 354.279p 10000.0u 354.28p 0 357.023p 0 357.024p 10000.0u 357.025p 0 359.153p 0 359.154p 10000.0u 359.155p 0 366.632p 0 366.633p 10000.0u 366.634p 0 368.657p 0 368.658p 10000.0u 368.659p 0 371.441p 0 371.442p 10000.0u 371.443p 0 381.434p 0 381.435p 10000.0u 381.436p 0 384.764p 0 384.765p 10000.0u 384.766p 0 391.49p 0 391.491p 10000.0u 391.492p 0 414.989p 0 414.99p 10000.0u 414.991p 0 418.016p 0 418.017p 10000.0u 418.018p 0 421.124p 0 421.125p 10000.0u 421.126p 0 425.42p 0 425.421p 10000.0u 425.422p 0 427.385p 0 427.386p 10000.0u 427.387p 0 436.625p 0 436.626p 10000.0u 436.627p 0 446.021p 0 446.022p 10000.0u 446.023p 0 447.716p 0 447.717p 10000.0u 447.718p 0 451.511p 0 451.512p 10000.0u 451.513p 0 472.235p 0 472.236p 10000.0u 472.237p 0 474.41p 0 474.411p 10000.0u 474.412p 0 486.032p 0 486.033p 10000.0u 486.034p 0 489.113p 0 489.114p 10000.0u 489.115p 0 500.948p 0 500.949p 10000.0u 500.95p 0 504.914p 0 504.915p 10000.0u 504.916p 0 505.643p 0 505.644p 10000.0u 505.645p 0 510.329p 0 510.33p 10000.0u 510.331p 0 523.511p 0 523.512p 10000.0u 523.513p 0 525.002p 0 525.003p 10000.0u 525.004p 0 525.281p 0 525.282p 10000.0u 525.283p 0 537.359p 0 537.36p 10000.0u 537.361p 0 545.99p 0 545.991p 10000.0u 545.992p 0 553.529p 0 553.53p 10000.0u 553.531p 0 556.352p 0 556.353p 10000.0u 556.354p 0 558.872p 0 558.873p 10000.0u 558.874p 0 589.982p 0 589.983p 10000.0u 589.984p 0 596.705p 0 596.706p 10000.0u 596.707p 0 603.854p 0 603.855p 10000.0u 603.856p 0 612.689p 0 612.69p 10000.0u 612.691p 0 624.674p 0 624.675p 10000.0u 624.676p 0 632.873p 0 632.874p 10000.0u 632.875p 0 639.356p 0 639.357p 10000.0u 639.358p 0 644.03p 0 644.031p 10000.0u 644.032p 0 652.235p 0 652.236p 10000.0u 652.237p 0 660.857p 0 660.858p 10000.0u 660.859p 0 661.163p 0 661.164p 10000.0u 661.165p 0 662.852p 0 662.853p 10000.0u 662.854p 0 664.964p 0 664.965p 10000.0u 664.966p 0 672.038p 0 672.039p 10000.0u 672.04p 0 679.508p 0 679.509p 10000.0u 679.51p 0 688.067p 0 688.068p 10000.0u 688.069p 0 693.977p 0 693.978p 10000.0u 693.979p 0 699.992p 0 699.993p 10000.0u 699.994p 0 720.644p 0 720.645p 10000.0u 720.646p 0 741.017p 0 741.018p 10000.0u 741.019p 0 743.579p 0 743.58p 10000.0u 743.581p 0 745.01p 0 745.011p 10000.0u 745.012p 0 755.372p 0 755.373p 10000.0u 755.374p 0 798.578p 0 798.579p 10000.0u 798.58p 0 836.366p 0 836.367p 10000.0u 836.368p 0 843.092p 0 843.093p 10000.0u 843.094p 0 860.255p 0 860.256p 10000.0u 860.257p 0 863.297p 0 863.298p 10000.0u 863.299p 0 869.234p 0 869.235p 10000.0u 869.236p 0 874.436p 0 874.437p 10000.0u 874.438p 0 876.773p 0 876.774p 10000.0u 876.775p 0 882.311p 0 882.312p 10000.0u 882.313p 0 883.124p 0 883.125p 10000.0u 883.126p 0 890.792p 0 890.793p 10000.0u 890.794p 0 908.837p 0 908.838p 10000.0u 908.839p 0 930.656p 0 930.657p 10000.0u 930.658p 0 949.307p 0 949.308p 10000.0u 949.309p 0 949.727p 0 949.728p 10000.0u 949.729p 0 961.031p 0 961.032p 10000.0u 961.033p 0 968.51p 0 968.511p 10000.0u 968.512p 0 991.43p 0 991.431p 10000.0u 991.432p 0 996.134p 0 996.135p 10000.0u 996.136p 0)
IIN17 0 18 pwl(0 0 31.757p 0 31.758p 10000.0u 31.759p 0 68.258p 0 68.259p 10000.0u 68.26p 0 71.285p 0 71.286p 10000.0u 71.287p 0 73.787p 0 73.788p 10000.0u 73.789p 0 87.542p 0 87.543p 10000.0u 87.544p 0 126.662p 0 126.663p 10000.0u 126.664p 0 134.981p 0 134.982p 10000.0u 134.983p 0 143.471p 0 143.472p 10000.0u 143.473p 0 151.973p 0 151.974p 10000.0u 151.975p 0 168.446p 0 168.447p 10000.0u 168.448p 0 173.345p 0 173.346p 10000.0u 173.347p 0 188.741p 0 188.742p 10000.0u 188.743p 0 203.864p 0 203.865p 10000.0u 203.866p 0 210.263p 0 210.264p 10000.0u 210.265p 0 215.48p 0 215.481p 10000.0u 215.482p 0 232.856p 0 232.857p 10000.0u 232.858p 0 234.824p 0 234.825p 10000.0u 234.826p 0 254.048p 0 254.049p 10000.0u 254.05p 0 257.384p 0 257.385p 10000.0u 257.386p 0 267.98p 0 267.981p 10000.0u 267.982p 0 282.887p 0 282.888p 10000.0u 282.889p 0 287.075p 0 287.076p 10000.0u 287.077p 0 292.391p 0 292.392p 10000.0u 292.393p 0 307.76p 0 307.761p 10000.0u 307.762p 0 308.279p 0 308.28p 10000.0u 308.281p 0 314.33p 0 314.331p 10000.0u 314.332p 0 330.632p 0 330.633p 10000.0u 330.634p 0 330.743p 0 330.744p 10000.0u 330.745p 0 336.62p 0 336.621p 10000.0u 336.622p 0 343.268p 0 343.269p 10000.0u 343.27p 0 371.399p 0 371.4p 10000.0u 371.401p 0 378.398p 0 378.399p 10000.0u 378.4p 0 392.432p 0 392.433p 10000.0u 392.434p 0 405.416p 0 405.417p 10000.0u 405.418p 0 423.473p 0 423.474p 10000.0u 423.475p 0 427.919p 0 427.92p 10000.0u 427.921p 0 441.914p 0 441.915p 10000.0u 441.916p 0 444.254p 0 444.255p 10000.0u 444.256p 0 446.672p 0 446.673p 10000.0u 446.674p 0 447.842p 0 447.843p 10000.0u 447.844p 0 461.609p 0 461.61p 10000.0u 461.611p 0 476.438p 0 476.439p 10000.0u 476.44p 0 483.86p 0 483.861p 10000.0u 483.862p 0 489.692p 0 489.693p 10000.0u 489.694p 0 494.9p 0 494.901p 10000.0u 494.902p 0 515.813p 0 515.814p 10000.0u 515.815p 0 518.381p 0 518.382p 10000.0u 518.383p 0 529.919p 0 529.92p 10000.0u 529.921p 0 548.801p 0 548.802p 10000.0u 548.803p 0 549.461p 0 549.462p 10000.0u 549.463p 0 552.458p 0 552.459p 10000.0u 552.46p 0 553.943p 0 553.944p 10000.0u 553.945p 0 563.945p 0 563.946p 10000.0u 563.947p 0 584.639p 0 584.64p 10000.0u 584.641p 0 594.506p 0 594.507p 10000.0u 594.508p 0 629.582p 0 629.583p 10000.0u 629.584p 0 641.861p 0 641.862p 10000.0u 641.863p 0 655.868p 0 655.869p 10000.0u 655.87p 0 656.963p 0 656.964p 10000.0u 656.965p 0 673.154p 0 673.155p 10000.0u 673.156p 0 685.067p 0 685.068p 10000.0u 685.069p 0 696.857p 0 696.858p 10000.0u 696.859p 0 706.394p 0 706.395p 10000.0u 706.396p 0 715.31p 0 715.311p 10000.0u 715.312p 0 728.246p 0 728.247p 10000.0u 728.248p 0 732.092p 0 732.093p 10000.0u 732.094p 0 732.311p 0 732.312p 10000.0u 732.313p 0 750.017p 0 750.018p 10000.0u 750.019p 0 754.418p 0 754.419p 10000.0u 754.42p 0 762.056p 0 762.057p 10000.0u 762.058p 0 770.591p 0 770.592p 10000.0u 770.593p 0 793.193p 0 793.194p 10000.0u 793.195p 0 793.997p 0 793.998p 10000.0u 793.999p 0 797.945p 0 797.946p 10000.0u 797.947p 0 802.022p 0 802.023p 10000.0u 802.024p 0 819.494p 0 819.495p 10000.0u 819.496p 0 821.315p 0 821.316p 10000.0u 821.317p 0 822.419p 0 822.42p 10000.0u 822.421p 0 841.952p 0 841.953p 10000.0u 841.954p 0 848.948p 0 848.949p 10000.0u 848.95p 0 855.449p 0 855.45p 10000.0u 855.451p 0 861.326p 0 861.327p 10000.0u 861.328p 0 865.643p 0 865.644p 10000.0u 865.645p 0 871.637p 0 871.638p 10000.0u 871.639p 0 891.347p 0 891.348p 10000.0u 891.349p 0 900.254p 0 900.255p 10000.0u 900.256p 0 918.827p 0 918.828p 10000.0u 918.829p 0 919.439p 0 919.44p 10000.0u 919.441p 0 926.78p 0 926.781p 10000.0u 926.782p 0 942.83p 0 942.831p 10000.0u 942.832p 0 952.469p 0 952.47p 10000.0u 952.471p 0 957.932p 0 957.933p 10000.0u 957.934p 0 983.594p 0 983.595p 10000.0u 983.596p 0)
IIN18 0 19 pwl(0 0 6.665p 0 6.666p 10000.0u 6.667p 0 11.987p 0 11.988p 10000.0u 11.989p 0 12.281p 0 12.282p 10000.0u 12.283p 0 14.024p 0 14.025p 10000.0u 14.026p 0 31.817p 0 31.818p 10000.0u 31.819p 0 41.45p 0 41.451p 10000.0u 41.452p 0 67.532p 0 67.533p 10000.0u 67.534p 0 72.761p 0 72.762p 10000.0u 72.763p 0 73.886p 0 73.887p 10000.0u 73.888p 0 97.55p 0 97.551p 10000.0u 97.552p 0 103.439p 0 103.44p 10000.0u 103.441p 0 112.835p 0 112.836p 10000.0u 112.837p 0 133.049p 0 133.05p 10000.0u 133.051p 0 133.853p 0 133.854p 10000.0u 133.855p 0 147.143p 0 147.144p 10000.0u 147.145p 0 153.854p 0 153.855p 10000.0u 153.856p 0 164.099p 0 164.1p 10000.0u 164.101p 0 166.799p 0 166.8p 10000.0u 166.801p 0 168.335p 0 168.336p 10000.0u 168.337p 0 180.938p 0 180.939p 10000.0u 180.94p 0 183.887p 0 183.888p 10000.0u 183.889p 0 188.783p 0 188.784p 10000.0u 188.785p 0 190.925p 0 190.926p 10000.0u 190.927p 0 204.098p 0 204.099p 10000.0u 204.1p 0 207.902p 0 207.903p 10000.0u 207.904p 0 212.786p 0 212.787p 10000.0u 212.788p 0 213.32p 0 213.321p 10000.0u 213.322p 0 233.615p 0 233.616p 10000.0u 233.617p 0 254.162p 0 254.163p 10000.0u 254.164p 0 259.676p 0 259.677p 10000.0u 259.678p 0 261.089p 0 261.09p 10000.0u 261.091p 0 263.936p 0 263.937p 10000.0u 263.938p 0 264.185p 0 264.186p 10000.0u 264.187p 0 271.376p 0 271.377p 10000.0u 271.378p 0 294.59p 0 294.591p 10000.0u 294.592p 0 297.971p 0 297.972p 10000.0u 297.973p 0 302.225p 0 302.226p 10000.0u 302.227p 0 315.368p 0 315.369p 10000.0u 315.37p 0 323.375p 0 323.376p 10000.0u 323.377p 0 328.601p 0 328.602p 10000.0u 328.603p 0 335.15p 0 335.151p 10000.0u 335.152p 0 348.188p 0 348.189p 10000.0u 348.19p 0 360.962p 0 360.963p 10000.0u 360.964p 0 370.823p 0 370.824p 10000.0u 370.825p 0 382.247p 0 382.248p 10000.0u 382.249p 0 384.908p 0 384.909p 10000.0u 384.91p 0 386.9p 0 386.901p 10000.0u 386.902p 0 392.171p 0 392.172p 10000.0u 392.173p 0 399.572p 0 399.573p 10000.0u 399.574p 0 404.333p 0 404.334p 10000.0u 404.335p 0 405.515p 0 405.516p 10000.0u 405.517p 0 431.051p 0 431.052p 10000.0u 431.053p 0 461.153p 0 461.154p 10000.0u 461.155p 0 472.184p 0 472.185p 10000.0u 472.186p 0 479.885p 0 479.886p 10000.0u 479.887p 0 485.39p 0 485.391p 10000.0u 485.392p 0 494.075p 0 494.076p 10000.0u 494.077p 0 498.188p 0 498.189p 10000.0u 498.19p 0 501.929p 0 501.93p 10000.0u 501.931p 0 503.771p 0 503.772p 10000.0u 503.773p 0 508.343p 0 508.344p 10000.0u 508.345p 0 509.06p 0 509.061p 10000.0u 509.062p 0 513.497p 0 513.498p 10000.0u 513.499p 0 540.911p 0 540.912p 10000.0u 540.913p 0 543.389p 0 543.39p 10000.0u 543.391p 0 548.975p 0 548.976p 10000.0u 548.977p 0 549.065p 0 549.066p 10000.0u 549.067p 0 566.372p 0 566.373p 10000.0u 566.374p 0 572.432p 0 572.433p 10000.0u 572.434p 0 573.872p 0 573.873p 10000.0u 573.874p 0 575.888p 0 575.889p 10000.0u 575.89p 0 583.13p 0 583.131p 10000.0u 583.132p 0 631.913p 0 631.914p 10000.0u 631.915p 0 649.943p 0 649.944p 10000.0u 649.945p 0 658.274p 0 658.275p 10000.0u 658.276p 0 665.912p 0 665.913p 10000.0u 665.914p 0 667.166p 0 667.167p 10000.0u 667.168p 0 675.584p 0 675.585p 10000.0u 675.586p 0 692.681p 0 692.682p 10000.0u 692.683p 0 694.652p 0 694.653p 10000.0u 694.654p 0 699.029p 0 699.03p 10000.0u 699.031p 0 701.033p 0 701.034p 10000.0u 701.035p 0 708.215p 0 708.216p 10000.0u 708.217p 0 723.755p 0 723.756p 10000.0u 723.757p 0 731.684p 0 731.685p 10000.0u 731.686p 0 735.407p 0 735.408p 10000.0u 735.409p 0 756.872p 0 756.873p 10000.0u 756.874p 0 768.917p 0 768.918p 10000.0u 768.919p 0 779.996p 0 779.997p 10000.0u 779.998p 0 783.167p 0 783.168p 10000.0u 783.169p 0 784.748p 0 784.749p 10000.0u 784.75p 0 790.955p 0 790.956p 10000.0u 790.957p 0 791.144p 0 791.145p 10000.0u 791.146p 0 792.596p 0 792.597p 10000.0u 792.598p 0 793.898p 0 793.899p 10000.0u 793.9p 0 803.57p 0 803.571p 10000.0u 803.572p 0 806.627p 0 806.628p 10000.0u 806.629p 0 808.79p 0 808.791p 10000.0u 808.792p 0 817.637p 0 817.638p 10000.0u 817.639p 0 844.4p 0 844.401p 10000.0u 844.402p 0 855.152p 0 855.153p 10000.0u 855.154p 0 861.557p 0 861.558p 10000.0u 861.559p 0 904.01p 0 904.011p 10000.0u 904.012p 0 921.128p 0 921.129p 10000.0u 921.13p 0 939.095p 0 939.096p 10000.0u 939.097p 0 940.607p 0 940.608p 10000.0u 940.609p 0 940.832p 0 940.833p 10000.0u 940.834p 0 954.113p 0 954.114p 10000.0u 954.115p 0 970.157p 0 970.158p 10000.0u 970.159p 0 976.328p 0 976.329p 10000.0u 976.33p 0 982.871p 0 982.872p 10000.0u 982.873p 0 995.216p 0 995.217p 10000.0u 995.218p 0 995.243p 0 995.244p 10000.0u 995.245p 0)
IIN19 0 20 pwl(0 0 15.845p 0 15.846p 10000.0u 15.847p 0 23.879p 0 23.88p 10000.0u 23.881p 0 37.307p 0 37.308p 10000.0u 37.309p 0 42.443p 0 42.444p 10000.0u 42.445p 0 46.547p 0 46.548p 10000.0u 46.549p 0 53.669p 0 53.67p 10000.0u 53.671p 0 66.308p 0 66.309p 10000.0u 66.31p 0 72.338p 0 72.339p 10000.0u 72.34p 0 73.448p 0 73.449p 10000.0u 73.45p 0 75.494p 0 75.495p 10000.0u 75.496p 0 82.694p 0 82.695p 10000.0u 82.696p 0 85.55p 0 85.551p 10000.0u 85.552p 0 110.606p 0 110.607p 10000.0u 110.608p 0 110.687p 0 110.688p 10000.0u 110.689p 0 121.745p 0 121.746p 10000.0u 121.747p 0 127.325p 0 127.326p 10000.0u 127.327p 0 129.287p 0 129.288p 10000.0u 129.289p 0 135.23p 0 135.231p 10000.0u 135.232p 0 143.843p 0 143.844p 10000.0u 143.845p 0 146.609p 0 146.61p 10000.0u 146.611p 0 163.694p 0 163.695p 10000.0u 163.696p 0 181.424p 0 181.425p 10000.0u 181.426p 0 183.602p 0 183.603p 10000.0u 183.604p 0 192.458p 0 192.459p 10000.0u 192.46p 0 203.408p 0 203.409p 10000.0u 203.41p 0 206.624p 0 206.625p 10000.0u 206.626p 0 210.881p 0 210.882p 10000.0u 210.883p 0 225.587p 0 225.588p 10000.0u 225.589p 0 242.423p 0 242.424p 10000.0u 242.425p 0 244.334p 0 244.335p 10000.0u 244.336p 0 254.474p 0 254.475p 10000.0u 254.476p 0 259.928p 0 259.929p 10000.0u 259.93p 0 268.265p 0 268.266p 10000.0u 268.267p 0 294.353p 0 294.354p 10000.0u 294.355p 0 306.041p 0 306.042p 10000.0u 306.043p 0 321.965p 0 321.966p 10000.0u 321.967p 0 325.049p 0 325.05p 10000.0u 325.051p 0 342.617p 0 342.618p 10000.0u 342.619p 0 353.003p 0 353.004p 10000.0u 353.005p 0 358.622p 0 358.623p 10000.0u 358.624p 0 370.313p 0 370.314p 10000.0u 370.315p 0 374.141p 0 374.142p 10000.0u 374.143p 0 382.139p 0 382.14p 10000.0u 382.141p 0 392.639p 0 392.64p 10000.0u 392.641p 0 416.42p 0 416.421p 10000.0u 416.422p 0 418.151p 0 418.152p 10000.0u 418.153p 0 423.914p 0 423.915p 10000.0u 423.916p 0 433.739p 0 433.74p 10000.0u 433.741p 0 440.438p 0 440.439p 10000.0u 440.44p 0 447.434p 0 447.435p 10000.0u 447.436p 0 456.95p 0 456.951p 10000.0u 456.952p 0 469.496p 0 469.497p 10000.0u 469.498p 0 474.116p 0 474.117p 10000.0u 474.118p 0 490.745p 0 490.746p 10000.0u 490.747p 0 522.509p 0 522.51p 10000.0u 522.511p 0 525.59p 0 525.591p 10000.0u 525.592p 0 530.858p 0 530.859p 10000.0u 530.86p 0 535.328p 0 535.329p 10000.0u 535.33p 0 543.704p 0 543.705p 10000.0u 543.706p 0 565.793p 0 565.794p 10000.0u 565.795p 0 570.989p 0 570.99p 10000.0u 570.991p 0 581.135p 0 581.136p 10000.0u 581.137p 0 603.164p 0 603.165p 10000.0u 603.166p 0 608.603p 0 608.604p 10000.0u 608.605p 0 624.767p 0 624.768p 10000.0u 624.769p 0 628.145p 0 628.146p 10000.0u 628.147p 0 629.759p 0 629.76p 10000.0u 629.761p 0 656.009p 0 656.01p 10000.0u 656.011p 0 657.365p 0 657.366p 10000.0u 657.367p 0 677.732p 0 677.733p 10000.0u 677.734p 0 681.404p 0 681.405p 10000.0u 681.406p 0 682.697p 0 682.698p 10000.0u 682.699p 0 688.124p 0 688.125p 10000.0u 688.126p 0 691.691p 0 691.692p 10000.0u 691.693p 0 700.367p 0 700.368p 10000.0u 700.369p 0 730.943p 0 730.944p 10000.0u 730.945p 0 765.809p 0 765.81p 10000.0u 765.811p 0 768.938p 0 768.939p 10000.0u 768.94p 0 786.038p 0 786.039p 10000.0u 786.04p 0 789.443p 0 789.444p 10000.0u 789.445p 0 807.803p 0 807.804p 10000.0u 807.805p 0 829.895p 0 829.896p 10000.0u 829.897p 0 840.302p 0 840.303p 10000.0u 840.304p 0 848.396p 0 848.397p 10000.0u 848.398p 0 900.665p 0 900.666p 10000.0u 900.667p 0 915.65p 0 915.651p 10000.0u 915.652p 0 919.202p 0 919.203p 10000.0u 919.204p 0 932.42p 0 932.421p 10000.0u 932.422p 0 932.528p 0 932.529p 10000.0u 932.53p 0 938.072p 0 938.073p 10000.0u 938.074p 0 944.036p 0 944.037p 10000.0u 944.038p 0 952.343p 0 952.344p 10000.0u 952.345p 0 964.205p 0 964.206p 10000.0u 964.207p 0 973.391p 0 973.392p 10000.0u 973.393p 0 980.825p 0 980.826p 10000.0u 980.827p 0 982.616p 0 982.617p 10000.0u 982.618p 0 983.174p 0 983.175p 10000.0u 983.176p 0 983.441p 0 983.442p 10000.0u 983.443p 0 997.016p 0 997.017p 10000.0u 997.018p 0)
IIN20 0 21 pwl(0 0 7.4p 0 7.401p 10000.0u 7.402p 0 34.679p 0 34.68p 10000.0u 34.681p 0 48.053p 0 48.054p 10000.0u 48.055p 0 50.579p 0 50.58p 10000.0u 50.581p 0 55.766p 0 55.767p 10000.0u 55.768p 0 72.176p 0 72.177p 10000.0u 72.178p 0 80.861p 0 80.862p 10000.0u 80.863p 0 110.306p 0 110.307p 10000.0u 110.308p 0 111.788p 0 111.789p 10000.0u 111.79p 0 128.279p 0 128.28p 10000.0u 128.281p 0 128.81p 0 128.811p 10000.0u 128.812p 0 130.964p 0 130.965p 10000.0u 130.966p 0 140.072p 0 140.073p 10000.0u 140.074p 0 147.905p 0 147.906p 10000.0u 147.907p 0 149.633p 0 149.634p 10000.0u 149.635p 0 164.627p 0 164.628p 10000.0u 164.629p 0 178.331p 0 178.332p 10000.0u 178.333p 0 181.019p 0 181.02p 10000.0u 181.021p 0 191.492p 0 191.493p 10000.0u 191.494p 0 203.333p 0 203.334p 10000.0u 203.335p 0 204.644p 0 204.645p 10000.0u 204.646p 0 213.074p 0 213.075p 10000.0u 213.076p 0 218.711p 0 218.712p 10000.0u 218.713p 0 227.489p 0 227.49p 10000.0u 227.491p 0 240.014p 0 240.015p 10000.0u 240.016p 0 247.952p 0 247.953p 10000.0u 247.954p 0 262.172p 0 262.173p 10000.0u 262.174p 0 262.763p 0 262.764p 10000.0u 262.765p 0 262.988p 0 262.989p 10000.0u 262.99p 0 266.072p 0 266.073p 10000.0u 266.074p 0 270.932p 0 270.933p 10000.0u 270.934p 0 275.87p 0 275.871p 10000.0u 275.872p 0 315.227p 0 315.228p 10000.0u 315.229p 0 317.369p 0 317.37p 10000.0u 317.371p 0 317.768p 0 317.769p 10000.0u 317.77p 0 319.331p 0 319.332p 10000.0u 319.333p 0 324.293p 0 324.294p 10000.0u 324.295p 0 336.47p 0 336.471p 10000.0u 336.472p 0 350.678p 0 350.679p 10000.0u 350.68p 0 354.32p 0 354.321p 10000.0u 354.322p 0 359.291p 0 359.292p 10000.0u 359.293p 0 361.025p 0 361.026p 10000.0u 361.027p 0 374.678p 0 374.679p 10000.0u 374.68p 0 418.133p 0 418.134p 10000.0u 418.135p 0 418.901p 0 418.902p 10000.0u 418.903p 0 431.348p 0 431.349p 10000.0u 431.35p 0 433.232p 0 433.233p 10000.0u 433.234p 0 442.805p 0 442.806p 10000.0u 442.807p 0 447.824p 0 447.825p 10000.0u 447.826p 0 453.833p 0 453.834p 10000.0u 453.835p 0 460.133p 0 460.134p 10000.0u 460.135p 0 460.595p 0 460.596p 10000.0u 460.597p 0 478.814p 0 478.815p 10000.0u 478.816p 0 490.187p 0 490.188p 10000.0u 490.189p 0 501.038p 0 501.039p 10000.0u 501.04p 0 505.34p 0 505.341p 10000.0u 505.342p 0 516.599p 0 516.6p 10000.0u 516.601p 0 520.817p 0 520.818p 10000.0u 520.819p 0 528.311p 0 528.312p 10000.0u 528.313p 0 538.706p 0 538.707p 10000.0u 538.708p 0 549.8p 0 549.801p 10000.0u 549.802p 0 559.361p 0 559.362p 10000.0u 559.363p 0 562.679p 0 562.68p 10000.0u 562.681p 0 564.656p 0 564.657p 10000.0u 564.658p 0 565.103p 0 565.104p 10000.0u 565.105p 0 576.569p 0 576.57p 10000.0u 576.571p 0 589.391p 0 589.392p 10000.0u 589.393p 0 591.758p 0 591.759p 10000.0u 591.76p 0 598.391p 0 598.392p 10000.0u 598.393p 0 603.527p 0 603.528p 10000.0u 603.529p 0 617.084p 0 617.085p 10000.0u 617.086p 0 637.316p 0 637.317p 10000.0u 637.318p 0 638.597p 0 638.598p 10000.0u 638.599p 0 641.978p 0 641.979p 10000.0u 641.98p 0 645.776p 0 645.777p 10000.0u 645.778p 0 646.022p 0 646.023p 10000.0u 646.024p 0 646.619p 0 646.62p 10000.0u 646.621p 0 654.626p 0 654.627p 10000.0u 654.628p 0 656.771p 0 656.772p 10000.0u 656.773p 0 660.212p 0 660.213p 10000.0u 660.214p 0 665.453p 0 665.454p 10000.0u 665.455p 0 680.816p 0 680.817p 10000.0u 680.818p 0 702.662p 0 702.663p 10000.0u 702.664p 0 709.091p 0 709.092p 10000.0u 709.093p 0 715.76p 0 715.761p 10000.0u 715.762p 0 721.163p 0 721.164p 10000.0u 721.165p 0 727.013p 0 727.014p 10000.0u 727.015p 0 732.596p 0 732.597p 10000.0u 732.598p 0 740.342p 0 740.343p 10000.0u 740.344p 0 753.464p 0 753.465p 10000.0u 753.466p 0 785.561p 0 785.562p 10000.0u 785.563p 0 785.651p 0 785.652p 10000.0u 785.653p 0 786.053p 0 786.054p 10000.0u 786.055p 0 790.274p 0 790.275p 10000.0u 790.276p 0 795.779p 0 795.78p 10000.0u 795.781p 0 796.283p 0 796.284p 10000.0u 796.285p 0 800.666p 0 800.667p 10000.0u 800.668p 0 810.071p 0 810.072p 10000.0u 810.073p 0 824.546p 0 824.547p 10000.0u 824.548p 0 849.476p 0 849.477p 10000.0u 849.478p 0 861.563p 0 861.564p 10000.0u 861.565p 0 871.346p 0 871.347p 10000.0u 871.348p 0 876.818p 0 876.819p 10000.0u 876.82p 0 879.047p 0 879.048p 10000.0u 879.049p 0 880.595p 0 880.596p 10000.0u 880.597p 0 883.037p 0 883.038p 10000.0u 883.039p 0 883.949p 0 883.95p 10000.0u 883.951p 0 890.42p 0 890.421p 10000.0u 890.422p 0 911.069p 0 911.07p 10000.0u 911.071p 0 917.612p 0 917.613p 10000.0u 917.614p 0 919.037p 0 919.038p 10000.0u 919.039p 0 931.1p 0 931.101p 10000.0u 931.102p 0 940.436p 0 940.437p 10000.0u 940.438p 0 965.315p 0 965.316p 10000.0u 965.317p 0 971.528p 0 971.529p 10000.0u 971.53p 0 976.247p 0 976.248p 10000.0u 976.249p 0 988.451p 0 988.452p 10000.0u 988.453p 0 989.639p 0 989.64p 10000.0u 989.641p 0)
IIN21 0 22 pwl(0 0 5.498p 0 5.499p 10000.0u 5.5p 0 17.771p 0 17.772p 10000.0u 17.773p 0 18.68p 0 18.681p 10000.0u 18.682p 0 22.439p 0 22.44p 10000.0u 22.441p 0 27.905p 0 27.906p 10000.0u 27.907p 0 36.149p 0 36.15p 10000.0u 36.151p 0 55.91p 0 55.911p 10000.0u 55.912p 0 60.173p 0 60.174p 10000.0u 60.175p 0 64.046p 0 64.047p 10000.0u 64.048p 0 69.578p 0 69.579p 10000.0u 69.58p 0 77.252p 0 77.253p 10000.0u 77.254p 0 79.487p 0 79.488p 10000.0u 79.489p 0 92.348p 0 92.349p 10000.0u 92.35p 0 98.642p 0 98.643p 10000.0u 98.644p 0 99.38p 0 99.381p 10000.0u 99.382p 0 123.299p 0 123.3p 10000.0u 123.301p 0 124.148p 0 124.149p 10000.0u 124.15p 0 135.35p 0 135.351p 10000.0u 135.352p 0 136.256p 0 136.257p 10000.0u 136.258p 0 146.135p 0 146.136p 10000.0u 146.137p 0 159.401p 0 159.402p 10000.0u 159.403p 0 173.351p 0 173.352p 10000.0u 173.353p 0 187.271p 0 187.272p 10000.0u 187.273p 0 187.952p 0 187.953p 10000.0u 187.954p 0 191.075p 0 191.076p 10000.0u 191.077p 0 192.407p 0 192.408p 10000.0u 192.409p 0 194.087p 0 194.088p 10000.0u 194.089p 0 194.864p 0 194.865p 10000.0u 194.866p 0 223.505p 0 223.506p 10000.0u 223.507p 0 228.398p 0 228.399p 10000.0u 228.4p 0 258.668p 0 258.669p 10000.0u 258.67p 0 260.606p 0 260.607p 10000.0u 260.608p 0 273.473p 0 273.474p 10000.0u 273.475p 0 285.788p 0 285.789p 10000.0u 285.79p 0 293.39p 0 293.391p 10000.0u 293.392p 0 310.433p 0 310.434p 10000.0u 310.435p 0 316.34p 0 316.341p 10000.0u 316.342p 0 319.685p 0 319.686p 10000.0u 319.687p 0 320.858p 0 320.859p 10000.0u 320.86p 0 322.421p 0 322.422p 10000.0u 322.423p 0 341.015p 0 341.016p 10000.0u 341.017p 0 363.815p 0 363.816p 10000.0u 363.817p 0 378.164p 0 378.165p 10000.0u 378.166p 0 378.269p 0 378.27p 10000.0u 378.271p 0 385.535p 0 385.536p 10000.0u 385.537p 0 387.26p 0 387.261p 10000.0u 387.262p 0 390.494p 0 390.495p 10000.0u 390.496p 0 399.734p 0 399.735p 10000.0u 399.736p 0 418.106p 0 418.107p 10000.0u 418.108p 0 421.583p 0 421.584p 10000.0u 421.585p 0 426.329p 0 426.33p 10000.0u 426.331p 0 443.543p 0 443.544p 10000.0u 443.545p 0 452.24p 0 452.241p 10000.0u 452.242p 0 453.596p 0 453.597p 10000.0u 453.598p 0 480.719p 0 480.72p 10000.0u 480.721p 0 483.137p 0 483.138p 10000.0u 483.139p 0 514.517p 0 514.518p 10000.0u 514.519p 0 519.203p 0 519.204p 10000.0u 519.205p 0 525.395p 0 525.396p 10000.0u 525.397p 0 526.847p 0 526.848p 10000.0u 526.849p 0 551.519p 0 551.52p 10000.0u 551.521p 0 557.294p 0 557.295p 10000.0u 557.296p 0 569.873p 0 569.874p 10000.0u 569.875p 0 600.374p 0 600.375p 10000.0u 600.376p 0 607.085p 0 607.086p 10000.0u 607.087p 0 607.973p 0 607.974p 10000.0u 607.975p 0 611.801p 0 611.802p 10000.0u 611.803p 0 622.334p 0 622.335p 10000.0u 622.336p 0 629.519p 0 629.52p 10000.0u 629.521p 0 637.892p 0 637.893p 10000.0u 637.894p 0 660.29p 0 660.291p 10000.0u 660.292p 0 690.968p 0 690.969p 10000.0u 690.97p 0 692.291p 0 692.292p 10000.0u 692.293p 0 709.127p 0 709.128p 10000.0u 709.129p 0 740.327p 0 740.328p 10000.0u 740.329p 0 740.915p 0 740.916p 10000.0u 740.917p 0 754.7p 0 754.701p 10000.0u 754.702p 0 787.772p 0 787.773p 10000.0u 787.774p 0 793.73p 0 793.731p 10000.0u 793.732p 0 804.767p 0 804.768p 10000.0u 804.769p 0 844.493p 0 844.494p 10000.0u 844.495p 0 847.64p 0 847.641p 10000.0u 847.642p 0 871.493p 0 871.494p 10000.0u 871.495p 0 902.57p 0 902.571p 10000.0u 902.572p 0 908.291p 0 908.292p 10000.0u 908.293p 0 911.531p 0 911.532p 10000.0u 911.533p 0 913.682p 0 913.683p 10000.0u 913.684p 0 923.561p 0 923.562p 10000.0u 923.563p 0 925.778p 0 925.779p 10000.0u 925.78p 0 935.435p 0 935.436p 10000.0u 935.437p 0 938.969p 0 938.97p 10000.0u 938.971p 0 949.535p 0 949.536p 10000.0u 949.537p 0 963.737p 0 963.738p 10000.0u 963.739p 0 989.795p 0 989.796p 10000.0u 989.797p 0 989.834p 0 989.835p 10000.0u 989.836p 0 998.948p 0 998.949p 10000.0u 998.95p 0)
IIN22 0 23 pwl(0 0 2.228p 0 2.229p 10000.0u 2.23p 0 8.657p 0 8.658p 10000.0u 8.659p 0 9.485p 0 9.486p 10000.0u 9.487p 0 42.767p 0 42.768p 10000.0u 42.769p 0 45.131p 0 45.132p 10000.0u 45.133p 0 88.298p 0 88.299p 10000.0u 88.3p 0 109.613p 0 109.614p 10000.0u 109.615p 0 119.222p 0 119.223p 10000.0u 119.224p 0 138.923p 0 138.924p 10000.0u 138.925p 0 147.497p 0 147.498p 10000.0u 147.499p 0 158.825p 0 158.826p 10000.0u 158.827p 0 169.049p 0 169.05p 10000.0u 169.051p 0 179.837p 0 179.838p 10000.0u 179.839p 0 182.042p 0 182.043p 10000.0u 182.044p 0 184.091p 0 184.092p 10000.0u 184.093p 0 186.887p 0 186.888p 10000.0u 186.889p 0 187.307p 0 187.308p 10000.0u 187.309p 0 215.951p 0 215.952p 10000.0u 215.953p 0 229.991p 0 229.992p 10000.0u 229.993p 0 250.742p 0 250.743p 10000.0u 250.744p 0 251.063p 0 251.064p 10000.0u 251.065p 0 254.642p 0 254.643p 10000.0u 254.644p 0 257.768p 0 257.769p 10000.0u 257.77p 0 269.348p 0 269.349p 10000.0u 269.35p 0 291.071p 0 291.072p 10000.0u 291.073p 0 299.642p 0 299.643p 10000.0u 299.644p 0 310.139p 0 310.14p 10000.0u 310.141p 0 310.946p 0 310.947p 10000.0u 310.948p 0 311.405p 0 311.406p 10000.0u 311.407p 0 341.699p 0 341.7p 10000.0u 341.701p 0 345.068p 0 345.069p 10000.0u 345.07p 0 348.458p 0 348.459p 10000.0u 348.46p 0 372.614p 0 372.615p 10000.0u 372.616p 0 373.874p 0 373.875p 10000.0u 373.876p 0 385.349p 0 385.35p 10000.0u 385.351p 0 387.77p 0 387.771p 10000.0u 387.772p 0 399.656p 0 399.657p 10000.0u 399.658p 0 405.824p 0 405.825p 10000.0u 405.826p 0 413.087p 0 413.088p 10000.0u 413.089p 0 429.404p 0 429.405p 10000.0u 429.406p 0 429.86p 0 429.861p 10000.0u 429.862p 0 437.87p 0 437.871p 10000.0u 437.872p 0 468.179p 0 468.18p 10000.0u 468.181p 0 471.125p 0 471.126p 10000.0u 471.127p 0 491.252p 0 491.253p 10000.0u 491.254p 0 495.809p 0 495.81p 10000.0u 495.811p 0 512.177p 0 512.178p 10000.0u 512.179p 0 534.701p 0 534.702p 10000.0u 534.703p 0 550.28p 0 550.281p 10000.0u 550.282p 0 551.531p 0 551.532p 10000.0u 551.533p 0 556.112p 0 556.113p 10000.0u 556.114p 0 557.177p 0 557.178p 10000.0u 557.179p 0 561.539p 0 561.54p 10000.0u 561.541p 0 562.307p 0 562.308p 10000.0u 562.309p 0 572.231p 0 572.232p 10000.0u 572.233p 0 586.283p 0 586.284p 10000.0u 586.285p 0 598.772p 0 598.773p 10000.0u 598.774p 0 599.645p 0 599.646p 10000.0u 599.647p 0 599.873p 0 599.874p 10000.0u 599.875p 0 612.644p 0 612.645p 10000.0u 612.646p 0 616.55p 0 616.551p 10000.0u 616.552p 0 642.092p 0 642.093p 10000.0u 642.094p 0 655.679p 0 655.68p 10000.0u 655.681p 0 668.207p 0 668.208p 10000.0u 668.209p 0 670.22p 0 670.221p 10000.0u 670.222p 0 671.681p 0 671.682p 10000.0u 671.683p 0 683.792p 0 683.793p 10000.0u 683.794p 0 691.331p 0 691.332p 10000.0u 691.333p 0 708.305p 0 708.306p 10000.0u 708.307p 0 741.452p 0 741.453p 10000.0u 741.454p 0 763.991p 0 763.992p 10000.0u 763.993p 0 785.645p 0 785.646p 10000.0u 785.647p 0 787.334p 0 787.335p 10000.0u 787.336p 0 792.785p 0 792.786p 10000.0u 792.787p 0 804.737p 0 804.738p 10000.0u 804.739p 0 815.612p 0 815.613p 10000.0u 815.614p 0 828.923p 0 828.924p 10000.0u 828.925p 0 867.359p 0 867.36p 10000.0u 867.361p 0 885.377p 0 885.378p 10000.0u 885.379p 0 915.803p 0 915.804p 10000.0u 915.805p 0 917.726p 0 917.727p 10000.0u 917.728p 0 922.631p 0 922.632p 10000.0u 922.633p 0 972.008p 0 972.009p 10000.0u 972.01p 0 976.757p 0 976.758p 10000.0u 976.759p 0 979.328p 0 979.329p 10000.0u 979.33p 0 980.0p 0 980.001p 10000.0u 980.002p 0)
IIN23 0 24 pwl(0 0 6.611p 0 6.612p 10000.0u 6.613p 0 23.576p 0 23.577p 10000.0u 23.578p 0 29.084p 0 29.085p 10000.0u 29.086p 0 35.465p 0 35.466p 10000.0u 35.467p 0 40.952p 0 40.953p 10000.0u 40.954p 0 60.617p 0 60.618p 10000.0u 60.619p 0 78.989p 0 78.99p 10000.0u 78.991p 0 80.249p 0 80.25p 10000.0u 80.251p 0 92.381p 0 92.382p 10000.0u 92.383p 0 96.194p 0 96.195p 10000.0u 96.196p 0 125.297p 0 125.298p 10000.0u 125.299p 0 136.715p 0 136.716p 10000.0u 136.717p 0 143.036p 0 143.037p 10000.0u 143.038p 0 146.159p 0 146.16p 10000.0u 146.161p 0 146.885p 0 146.886p 10000.0u 146.887p 0 159.5p 0 159.501p 10000.0u 159.502p 0 164.9p 0 164.901p 10000.0u 164.902p 0 170.708p 0 170.709p 10000.0u 170.71p 0 172.289p 0 172.29p 10000.0u 172.291p 0 178.979p 0 178.98p 10000.0u 178.981p 0 182.225p 0 182.226p 10000.0u 182.227p 0 193.919p 0 193.92p 10000.0u 193.921p 0 211.667p 0 211.668p 10000.0u 211.669p 0 231.917p 0 231.918p 10000.0u 231.919p 0 241.892p 0 241.893p 10000.0u 241.894p 0 242.783p 0 242.784p 10000.0u 242.785p 0 243.929p 0 243.93p 10000.0u 243.931p 0 250.511p 0 250.512p 10000.0u 250.513p 0 254.84p 0 254.841p 10000.0u 254.842p 0 267.362p 0 267.363p 10000.0u 267.364p 0 282.104p 0 282.105p 10000.0u 282.106p 0 295.298p 0 295.299p 10000.0u 295.3p 0 302.897p 0 302.898p 10000.0u 302.899p 0 313.685p 0 313.686p 10000.0u 313.687p 0 320.153p 0 320.154p 10000.0u 320.155p 0 329.978p 0 329.979p 10000.0u 329.98p 0 331.118p 0 331.119p 10000.0u 331.12p 0 356.942p 0 356.943p 10000.0u 356.944p 0 357.623p 0 357.624p 10000.0u 357.625p 0 365.828p 0 365.829p 10000.0u 365.83p 0 366.986p 0 366.987p 10000.0u 366.988p 0 377.984p 0 377.985p 10000.0u 377.986p 0 378.308p 0 378.309p 10000.0u 378.31p 0 392.42p 0 392.421p 10000.0u 392.422p 0 408.794p 0 408.795p 10000.0u 408.796p 0 416.426p 0 416.427p 10000.0u 416.428p 0 424.352p 0 424.353p 10000.0u 424.354p 0 427.199p 0 427.2p 10000.0u 427.201p 0 438.614p 0 438.615p 10000.0u 438.616p 0 444.818p 0 444.819p 10000.0u 444.82p 0 453.173p 0 453.174p 10000.0u 453.175p 0 455.756p 0 455.757p 10000.0u 455.758p 0 493.913p 0 493.914p 10000.0u 493.915p 0 495.632p 0 495.633p 10000.0u 495.634p 0 523.574p 0 523.575p 10000.0u 523.576p 0 526.487p 0 526.488p 10000.0u 526.489p 0 536.759p 0 536.76p 10000.0u 536.761p 0 542.102p 0 542.103p 10000.0u 542.104p 0 542.915p 0 542.916p 10000.0u 542.917p 0 547.151p 0 547.152p 10000.0u 547.153p 0 561.353p 0 561.354p 10000.0u 561.355p 0 566.576p 0 566.577p 10000.0u 566.578p 0 568.223p 0 568.224p 10000.0u 568.225p 0 586.76p 0 586.761p 10000.0u 586.762p 0 620.735p 0 620.736p 10000.0u 620.737p 0 623.927p 0 623.928p 10000.0u 623.929p 0 626.882p 0 626.883p 10000.0u 626.884p 0 630.161p 0 630.162p 10000.0u 630.163p 0 640.625p 0 640.626p 10000.0u 640.627p 0 647.957p 0 647.958p 10000.0u 647.959p 0 651.629p 0 651.63p 10000.0u 651.631p 0 656.489p 0 656.49p 10000.0u 656.491p 0 661.058p 0 661.059p 10000.0u 661.06p 0 697.379p 0 697.38p 10000.0u 697.381p 0 716.486p 0 716.487p 10000.0u 716.488p 0 718.025p 0 718.026p 10000.0u 718.027p 0 763.829p 0 763.83p 10000.0u 763.831p 0 764.375p 0 764.376p 10000.0u 764.377p 0 772.088p 0 772.089p 10000.0u 772.09p 0 777.401p 0 777.402p 10000.0u 777.403p 0 803.549p 0 803.55p 10000.0u 803.551p 0 809.057p 0 809.058p 10000.0u 809.059p 0 817.448p 0 817.449p 10000.0u 817.45p 0 827.126p 0 827.127p 10000.0u 827.128p 0 827.99p 0 827.991p 10000.0u 827.992p 0 836.966p 0 836.967p 10000.0u 836.968p 0 837.305p 0 837.306p 10000.0u 837.307p 0 839.651p 0 839.652p 10000.0u 839.653p 0 844.901p 0 844.902p 10000.0u 844.903p 0 866.798p 0 866.799p 10000.0u 866.8p 0 868.904p 0 868.905p 10000.0u 868.906p 0 883.553p 0 883.554p 10000.0u 883.555p 0 886.583p 0 886.584p 10000.0u 886.585p 0 887.432p 0 887.433p 10000.0u 887.434p 0 888.569p 0 888.57p 10000.0u 888.571p 0 891.68p 0 891.681p 10000.0u 891.682p 0 914.993p 0 914.994p 10000.0u 914.995p 0 946.223p 0 946.224p 10000.0u 946.225p 0 946.454p 0 946.455p 10000.0u 946.456p 0 953.543p 0 953.544p 10000.0u 953.545p 0 956.552p 0 956.553p 10000.0u 956.554p 0 961.565p 0 961.566p 10000.0u 961.567p 0 962.87p 0 962.871p 10000.0u 962.872p 0)
IIN24 0 25 pwl(0 0 18.269p 0 18.27p 10000.0u 18.271p 0 20.765p 0 20.766p 10000.0u 20.767p 0 58.73p 0 58.731p 10000.0u 58.732p 0 76.868p 0 76.869p 10000.0u 76.87p 0 85.61p 0 85.611p 10000.0u 85.612p 0 109.604p 0 109.605p 10000.0u 109.606p 0 129.176p 0 129.177p 10000.0u 129.178p 0 152.534p 0 152.535p 10000.0u 152.536p 0 188.906p 0 188.907p 10000.0u 188.908p 0 196.844p 0 196.845p 10000.0u 196.846p 0 200.456p 0 200.457p 10000.0u 200.458p 0 208.4p 0 208.401p 10000.0u 208.402p 0 217.199p 0 217.2p 10000.0u 217.201p 0 218.27p 0 218.271p 10000.0u 218.272p 0 221.204p 0 221.205p 10000.0u 221.206p 0 221.282p 0 221.283p 10000.0u 221.284p 0 231.908p 0 231.909p 10000.0u 231.91p 0 233.393p 0 233.394p 10000.0u 233.395p 0 235.196p 0 235.197p 10000.0u 235.198p 0 236.735p 0 236.736p 10000.0u 236.737p 0 237.098p 0 237.099p 10000.0u 237.1p 0 253.73p 0 253.731p 10000.0u 253.732p 0 260.039p 0 260.04p 10000.0u 260.041p 0 273.785p 0 273.786p 10000.0u 273.787p 0 284.384p 0 284.385p 10000.0u 284.386p 0 285.596p 0 285.597p 10000.0u 285.598p 0 294.515p 0 294.516p 10000.0u 294.517p 0 318.32p 0 318.321p 10000.0u 318.322p 0 318.563p 0 318.564p 10000.0u 318.565p 0 334.079p 0 334.08p 10000.0u 334.081p 0 335.813p 0 335.814p 10000.0u 335.815p 0 340.004p 0 340.005p 10000.0u 340.006p 0 348.449p 0 348.45p 10000.0u 348.451p 0 354.152p 0 354.153p 10000.0u 354.154p 0 355.163p 0 355.164p 10000.0u 355.165p 0 361.331p 0 361.332p 10000.0u 361.333p 0 380.456p 0 380.457p 10000.0u 380.458p 0 392.285p 0 392.286p 10000.0u 392.287p 0 394.787p 0 394.788p 10000.0u 394.789p 0 395.081p 0 395.082p 10000.0u 395.083p 0 396.872p 0 396.873p 10000.0u 396.874p 0 411.809p 0 411.81p 10000.0u 411.811p 0 435.449p 0 435.45p 10000.0u 435.451p 0 456.98p 0 456.981p 10000.0u 456.982p 0 460.196p 0 460.197p 10000.0u 460.198p 0 462.674p 0 462.675p 10000.0u 462.676p 0 464.54p 0 464.541p 10000.0u 464.542p 0 480.128p 0 480.129p 10000.0u 480.13p 0 481.022p 0 481.023p 10000.0u 481.024p 0 499.523p 0 499.524p 10000.0u 499.525p 0 511.262p 0 511.263p 10000.0u 511.264p 0 512.087p 0 512.088p 10000.0u 512.089p 0 516.776p 0 516.777p 10000.0u 516.778p 0 519.899p 0 519.9p 10000.0u 519.901p 0 523.592p 0 523.593p 10000.0u 523.594p 0 531.416p 0 531.417p 10000.0u 531.418p 0 541.838p 0 541.839p 10000.0u 541.84p 0 548.357p 0 548.358p 10000.0u 548.359p 0 554.354p 0 554.355p 10000.0u 554.356p 0 554.687p 0 554.688p 10000.0u 554.689p 0 574.097p 0 574.098p 10000.0u 574.099p 0 613.028p 0 613.029p 10000.0u 613.03p 0 623.135p 0 623.136p 10000.0u 623.137p 0 635.522p 0 635.523p 10000.0u 635.524p 0 643.082p 0 643.083p 10000.0u 643.084p 0 644.351p 0 644.352p 10000.0u 644.353p 0 646.946p 0 646.947p 10000.0u 646.948p 0 659.117p 0 659.118p 10000.0u 659.119p 0 679.883p 0 679.884p 10000.0u 679.885p 0 686.924p 0 686.925p 10000.0u 686.926p 0 704.96p 0 704.961p 10000.0u 704.962p 0 710.168p 0 710.169p 10000.0u 710.17p 0 727.733p 0 727.734p 10000.0u 727.735p 0 735.284p 0 735.285p 10000.0u 735.286p 0 736.025p 0 736.026p 10000.0u 736.027p 0 740.339p 0 740.34p 10000.0u 740.341p 0 755.114p 0 755.115p 10000.0u 755.116p 0 756.059p 0 756.06p 10000.0u 756.061p 0 769.679p 0 769.68p 10000.0u 769.681p 0 776.048p 0 776.049p 10000.0u 776.05p 0 776.744p 0 776.745p 10000.0u 776.746p 0 788.876p 0 788.877p 10000.0u 788.878p 0 789.197p 0 789.198p 10000.0u 789.199p 0 790.844p 0 790.845p 10000.0u 790.846p 0 793.04p 0 793.041p 10000.0u 793.042p 0 813.377p 0 813.378p 10000.0u 813.379p 0 814.892p 0 814.893p 10000.0u 814.894p 0 821.132p 0 821.133p 10000.0u 821.134p 0 821.819p 0 821.82p 10000.0u 821.821p 0 845.603p 0 845.604p 10000.0u 845.605p 0 863.567p 0 863.568p 10000.0u 863.569p 0 865.184p 0 865.185p 10000.0u 865.186p 0 876.335p 0 876.336p 10000.0u 876.337p 0 894.128p 0 894.129p 10000.0u 894.13p 0 894.692p 0 894.693p 10000.0u 894.694p 0 900.236p 0 900.237p 10000.0u 900.238p 0 900.764p 0 900.765p 10000.0u 900.766p 0 903.467p 0 903.468p 10000.0u 903.469p 0 904.601p 0 904.602p 10000.0u 904.603p 0 923.423p 0 923.424p 10000.0u 923.425p 0 938.27p 0 938.271p 10000.0u 938.272p 0 944.075p 0 944.076p 10000.0u 944.077p 0 986.693p 0 986.694p 10000.0u 986.695p 0 996.383p 0 996.384p 10000.0u 996.385p 0)
IIN25 0 26 pwl(0 0 9.728p 0 9.729p 10000.0u 9.73p 0 15.167p 0 15.168p 10000.0u 15.169p 0 29.672p 0 29.673p 10000.0u 29.674p 0 43.859p 0 43.86p 10000.0u 43.861p 0 48.563p 0 48.564p 10000.0u 48.565p 0 53.531p 0 53.532p 10000.0u 53.533p 0 66.299p 0 66.3p 10000.0u 66.301p 0 72.293p 0 72.294p 10000.0u 72.295p 0 85.733p 0 85.734p 10000.0u 85.735p 0 91.094p 0 91.095p 10000.0u 91.096p 0 91.958p 0 91.959p 10000.0u 91.96p 0 102.803p 0 102.804p 10000.0u 102.805p 0 108.569p 0 108.57p 10000.0u 108.571p 0 109.286p 0 109.287p 10000.0u 109.288p 0 129.809p 0 129.81p 10000.0u 129.811p 0 142.787p 0 142.788p 10000.0u 142.789p 0 146.633p 0 146.634p 10000.0u 146.635p 0 160.331p 0 160.332p 10000.0u 160.333p 0 169.853p 0 169.854p 10000.0u 169.855p 0 187.511p 0 187.512p 10000.0u 187.513p 0 188.954p 0 188.955p 10000.0u 188.956p 0 189.899p 0 189.9p 10000.0u 189.901p 0 190.982p 0 190.983p 10000.0u 190.984p 0 203.954p 0 203.955p 10000.0u 203.956p 0 207.029p 0 207.03p 10000.0u 207.031p 0 209.369p 0 209.37p 10000.0u 209.371p 0 211.865p 0 211.866p 10000.0u 211.867p 0 224.417p 0 224.418p 10000.0u 224.419p 0 227.027p 0 227.028p 10000.0u 227.029p 0 262.811p 0 262.812p 10000.0u 262.813p 0 268.379p 0 268.38p 10000.0u 268.381p 0 273.989p 0 273.99p 10000.0u 273.991p 0 278.747p 0 278.748p 10000.0u 278.749p 0 293.744p 0 293.745p 10000.0u 293.746p 0 309.995p 0 309.996p 10000.0u 309.997p 0 312.353p 0 312.354p 10000.0u 312.355p 0 323.723p 0 323.724p 10000.0u 323.725p 0 323.738p 0 323.739p 10000.0u 323.74p 0 328.481p 0 328.482p 10000.0u 328.483p 0 337.265p 0 337.266p 10000.0u 337.267p 0 345.674p 0 345.675p 10000.0u 345.676p 0 348.002p 0 348.003p 10000.0u 348.004p 0 355.085p 0 355.086p 10000.0u 355.087p 0 356.378p 0 356.379p 10000.0u 356.38p 0 362.717p 0 362.718p 10000.0u 362.719p 0 371.387p 0 371.388p 10000.0u 371.389p 0 381.533p 0 381.534p 10000.0u 381.535p 0 389.996p 0 389.997p 10000.0u 389.998p 0 396.929p 0 396.93p 10000.0u 396.931p 0 401.156p 0 401.157p 10000.0u 401.158p 0 418.064p 0 418.065p 10000.0u 418.066p 0 423.383p 0 423.384p 10000.0u 423.385p 0 429.383p 0 429.384p 10000.0u 429.385p 0 435.104p 0 435.105p 10000.0u 435.106p 0 437.837p 0 437.838p 10000.0u 437.839p 0 440.81p 0 440.811p 10000.0u 440.812p 0 479.858p 0 479.859p 10000.0u 479.86p 0 496.244p 0 496.245p 10000.0u 496.246p 0 506.18p 0 506.181p 10000.0u 506.182p 0 514.766p 0 514.767p 10000.0u 514.768p 0 519.521p 0 519.522p 10000.0u 519.523p 0 523.649p 0 523.65p 10000.0u 523.651p 0 525.164p 0 525.165p 10000.0u 525.166p 0 547.652p 0 547.653p 10000.0u 547.654p 0 554.111p 0 554.112p 10000.0u 554.113p 0 564.395p 0 564.396p 10000.0u 564.397p 0 576.164p 0 576.165p 10000.0u 576.166p 0 577.274p 0 577.275p 10000.0u 577.276p 0 589.253p 0 589.254p 10000.0u 589.255p 0 603.395p 0 603.396p 10000.0u 603.397p 0 618.452p 0 618.453p 10000.0u 618.454p 0 624.665p 0 624.666p 10000.0u 624.667p 0 628.055p 0 628.056p 10000.0u 628.057p 0 644.72p 0 644.721p 10000.0u 644.722p 0 652.118p 0 652.119p 10000.0u 652.12p 0 664.616p 0 664.617p 10000.0u 664.618p 0 666.56p 0 666.561p 10000.0u 666.562p 0 666.947p 0 666.948p 10000.0u 666.949p 0 672.818p 0 672.819p 10000.0u 672.82p 0 687.494p 0 687.495p 10000.0u 687.496p 0 687.749p 0 687.75p 10000.0u 687.751p 0 702.56p 0 702.561p 10000.0u 702.562p 0 716.675p 0 716.676p 10000.0u 716.677p 0 724.472p 0 724.473p 10000.0u 724.474p 0 726.377p 0 726.378p 10000.0u 726.379p 0 727.232p 0 727.233p 10000.0u 727.234p 0 731.801p 0 731.802p 10000.0u 731.803p 0 738.533p 0 738.534p 10000.0u 738.535p 0 752.96p 0 752.961p 10000.0u 752.962p 0 772.943p 0 772.944p 10000.0u 772.945p 0 778.112p 0 778.113p 10000.0u 778.114p 0 780.56p 0 780.561p 10000.0u 780.562p 0 788.342p 0 788.343p 10000.0u 788.344p 0 791.537p 0 791.538p 10000.0u 791.539p 0 799.142p 0 799.143p 10000.0u 799.144p 0 813.404p 0 813.405p 10000.0u 813.406p 0 814.589p 0 814.59p 10000.0u 814.591p 0 817.013p 0 817.014p 10000.0u 817.015p 0 833.006p 0 833.007p 10000.0u 833.008p 0 849.53p 0 849.531p 10000.0u 849.532p 0 850.685p 0 850.686p 10000.0u 850.687p 0 870.95p 0 870.951p 10000.0u 870.952p 0 877.076p 0 877.077p 10000.0u 877.078p 0 878.132p 0 878.133p 10000.0u 878.134p 0 884.705p 0 884.706p 10000.0u 884.707p 0 893.885p 0 893.886p 10000.0u 893.887p 0 916.388p 0 916.389p 10000.0u 916.39p 0 929.177p 0 929.178p 10000.0u 929.179p 0 935.042p 0 935.043p 10000.0u 935.044p 0 935.783p 0 935.784p 10000.0u 935.785p 0 949.988p 0 949.989p 10000.0u 949.99p 0 953.843p 0 953.844p 10000.0u 953.845p 0 965.186p 0 965.187p 10000.0u 965.188p 0 965.531p 0 965.532p 10000.0u 965.533p 0 981.176p 0 981.177p 10000.0u 981.178p 0 981.536p 0 981.537p 10000.0u 981.538p 0 983.333p 0 983.334p 10000.0u 983.335p 0 986.075p 0 986.076p 10000.0u 986.077p 0 991.151p 0 991.152p 10000.0u 991.153p 0)
IIN26 0 27 pwl(0 0 2.837p 0 2.838p 10000.0u 2.839p 0 5.297p 0 5.298p 10000.0u 5.299p 0 6.833p 0 6.834p 10000.0u 6.835p 0 8.594p 0 8.595p 10000.0u 8.596p 0 28.022p 0 28.023p 10000.0u 28.024p 0 39.272p 0 39.273p 10000.0u 39.274p 0 56.387p 0 56.388p 10000.0u 56.389p 0 60.098p 0 60.099p 10000.0u 60.1p 0 83.18p 0 83.181p 10000.0u 83.182p 0 86.057p 0 86.058p 10000.0u 86.059p 0 93.773p 0 93.774p 10000.0u 93.775p 0 102.65p 0 102.651p 10000.0u 102.652p 0 115.427p 0 115.428p 10000.0u 115.429p 0 121.547p 0 121.548p 10000.0u 121.549p 0 129.386p 0 129.387p 10000.0u 129.388p 0 148.637p 0 148.638p 10000.0u 148.639p 0 159.824p 0 159.825p 10000.0u 159.826p 0 160.202p 0 160.203p 10000.0u 160.204p 0 160.928p 0 160.929p 10000.0u 160.93p 0 164.207p 0 164.208p 10000.0u 164.209p 0 201.155p 0 201.156p 10000.0u 201.157p 0 212.075p 0 212.076p 10000.0u 212.077p 0 273.434p 0 273.435p 10000.0u 273.436p 0 297.773p 0 297.774p 10000.0u 297.775p 0 311.129p 0 311.13p 10000.0u 311.131p 0 330.125p 0 330.126p 10000.0u 330.127p 0 334.664p 0 334.665p 10000.0u 334.666p 0 338.201p 0 338.202p 10000.0u 338.203p 0 357.329p 0 357.33p 10000.0u 357.331p 0 364.685p 0 364.686p 10000.0u 364.687p 0 375.287p 0 375.288p 10000.0u 375.289p 0 386.807p 0 386.808p 10000.0u 386.809p 0 388.292p 0 388.293p 10000.0u 388.294p 0 399.731p 0 399.732p 10000.0u 399.733p 0 401.981p 0 401.982p 10000.0u 401.983p 0 403.724p 0 403.725p 10000.0u 403.726p 0 420.311p 0 420.312p 10000.0u 420.313p 0 427.181p 0 427.182p 10000.0u 427.183p 0 438.704p 0 438.705p 10000.0u 438.706p 0 441.662p 0 441.663p 10000.0u 441.664p 0 454.814p 0 454.815p 10000.0u 454.816p 0 457.499p 0 457.5p 10000.0u 457.501p 0 471.278p 0 471.279p 10000.0u 471.28p 0 501.167p 0 501.168p 10000.0u 501.169p 0 502.745p 0 502.746p 10000.0u 502.747p 0 506.615p 0 506.616p 10000.0u 506.617p 0 509.885p 0 509.886p 10000.0u 509.887p 0 529.652p 0 529.653p 10000.0u 529.654p 0 541.115p 0 541.116p 10000.0u 541.117p 0 548.198p 0 548.199p 10000.0u 548.2p 0 560.582p 0 560.583p 10000.0u 560.584p 0 564.854p 0 564.855p 10000.0u 564.856p 0 565.838p 0 565.839p 10000.0u 565.84p 0 569.327p 0 569.328p 10000.0u 569.329p 0 570.44p 0 570.441p 10000.0u 570.442p 0 632.468p 0 632.469p 10000.0u 632.47p 0 672.809p 0 672.81p 10000.0u 672.811p 0 683.351p 0 683.352p 10000.0u 683.353p 0 685.775p 0 685.776p 10000.0u 685.777p 0 688.571p 0 688.572p 10000.0u 688.573p 0 703.202p 0 703.203p 10000.0u 703.204p 0 710.45p 0 710.451p 10000.0u 710.452p 0 718.118p 0 718.119p 10000.0u 718.12p 0 738.929p 0 738.93p 10000.0u 738.931p 0 741.233p 0 741.234p 10000.0u 741.235p 0 751.247p 0 751.248p 10000.0u 751.249p 0 761.846p 0 761.847p 10000.0u 761.848p 0 769.535p 0 769.536p 10000.0u 769.537p 0 771.308p 0 771.309p 10000.0u 771.31p 0 788.243p 0 788.244p 10000.0u 788.245p 0 791.417p 0 791.418p 10000.0u 791.419p 0 791.678p 0 791.679p 10000.0u 791.68p 0 838.241p 0 838.242p 10000.0u 838.243p 0 842.435p 0 842.436p 10000.0u 842.437p 0 860.792p 0 860.793p 10000.0u 860.794p 0 869.219p 0 869.22p 10000.0u 869.221p 0 873.731p 0 873.732p 10000.0u 873.733p 0 883.373p 0 883.374p 10000.0u 883.375p 0 909.656p 0 909.657p 10000.0u 909.658p 0 938.624p 0 938.625p 10000.0u 938.626p 0 946.922p 0 946.923p 10000.0u 946.924p 0 968.318p 0 968.319p 10000.0u 968.32p 0 994.064p 0 994.065p 10000.0u 994.066p 0 998.849p 0 998.85p 10000.0u 998.851p 0)
IIN27 0 28 pwl(0 0 30.647p 0 30.648p 10000.0u 30.649p 0 43.91p 0 43.911p 10000.0u 43.912p 0 54.296p 0 54.297p 10000.0u 54.298p 0 79.331p 0 79.332p 10000.0u 79.333p 0 87.878p 0 87.879p 10000.0u 87.88p 0 89.279p 0 89.28p 10000.0u 89.281p 0 116.375p 0 116.376p 10000.0u 116.377p 0 117.557p 0 117.558p 10000.0u 117.559p 0 129.266p 0 129.267p 10000.0u 129.268p 0 139.703p 0 139.704p 10000.0u 139.705p 0 144.911p 0 144.912p 10000.0u 144.913p 0 151.67p 0 151.671p 10000.0u 151.672p 0 157.865p 0 157.866p 10000.0u 157.867p 0 163.283p 0 163.284p 10000.0u 163.285p 0 170.474p 0 170.475p 10000.0u 170.476p 0 173.519p 0 173.52p 10000.0u 173.521p 0 173.927p 0 173.928p 10000.0u 173.929p 0 174.995p 0 174.996p 10000.0u 174.997p 0 179.297p 0 179.298p 10000.0u 179.299p 0 195.989p 0 195.99p 10000.0u 195.991p 0 199.079p 0 199.08p 10000.0u 199.081p 0 208.916p 0 208.917p 10000.0u 208.918p 0 211.04p 0 211.041p 10000.0u 211.042p 0 215.942p 0 215.943p 10000.0u 215.944p 0 217.343p 0 217.344p 10000.0u 217.345p 0 225.938p 0 225.939p 10000.0u 225.94p 0 243.077p 0 243.078p 10000.0u 243.079p 0 246.362p 0 246.363p 10000.0u 246.364p 0 251.105p 0 251.106p 10000.0u 251.107p 0 257.801p 0 257.802p 10000.0u 257.803p 0 265.418p 0 265.419p 10000.0u 265.42p 0 287.237p 0 287.238p 10000.0u 287.239p 0 293.804p 0 293.805p 10000.0u 293.806p 0 294.221p 0 294.222p 10000.0u 294.223p 0 305.546p 0 305.547p 10000.0u 305.548p 0 307.625p 0 307.626p 10000.0u 307.627p 0 342.257p 0 342.258p 10000.0u 342.259p 0 351.584p 0 351.585p 10000.0u 351.586p 0 353.747p 0 353.748p 10000.0u 353.749p 0 354.674p 0 354.675p 10000.0u 354.676p 0 355.709p 0 355.71p 10000.0u 355.711p 0 355.871p 0 355.872p 10000.0u 355.873p 0 362.858p 0 362.859p 10000.0u 362.86p 0 376.631p 0 376.632p 10000.0u 376.633p 0 376.763p 0 376.764p 10000.0u 376.765p 0 384.341p 0 384.342p 10000.0u 384.343p 0 391.22p 0 391.221p 10000.0u 391.222p 0 391.421p 0 391.422p 10000.0u 391.423p 0 392.183p 0 392.184p 10000.0u 392.185p 0 394.244p 0 394.245p 10000.0u 394.246p 0 404.957p 0 404.958p 10000.0u 404.959p 0 417.737p 0 417.738p 10000.0u 417.739p 0 423.143p 0 423.144p 10000.0u 423.145p 0 432.716p 0 432.717p 10000.0u 432.718p 0 433.112p 0 433.113p 10000.0u 433.114p 0 449.156p 0 449.157p 10000.0u 449.158p 0 473.972p 0 473.973p 10000.0u 473.974p 0 478.202p 0 478.203p 10000.0u 478.204p 0 478.382p 0 478.383p 10000.0u 478.384p 0 485.75p 0 485.751p 10000.0u 485.752p 0 486.152p 0 486.153p 10000.0u 486.154p 0 507.497p 0 507.498p 10000.0u 507.499p 0 507.776p 0 507.777p 10000.0u 507.778p 0 521.348p 0 521.349p 10000.0u 521.35p 0 522.347p 0 522.348p 10000.0u 522.349p 0 522.881p 0 522.882p 10000.0u 522.883p 0 537.623p 0 537.624p 10000.0u 537.625p 0 539.381p 0 539.382p 10000.0u 539.383p 0 554.288p 0 554.289p 10000.0u 554.29p 0 556.688p 0 556.689p 10000.0u 556.69p 0 558.632p 0 558.633p 10000.0u 558.634p 0 574.499p 0 574.5p 10000.0u 574.501p 0 576.11p 0 576.111p 10000.0u 576.112p 0 595.025p 0 595.026p 10000.0u 595.027p 0 597.776p 0 597.777p 10000.0u 597.778p 0 601.151p 0 601.152p 10000.0u 601.153p 0 607.325p 0 607.326p 10000.0u 607.327p 0 610.448p 0 610.449p 10000.0u 610.45p 0 618.191p 0 618.192p 10000.0u 618.193p 0 618.314p 0 618.315p 10000.0u 618.316p 0 623.678p 0 623.679p 10000.0u 623.68p 0 632.552p 0 632.553p 10000.0u 632.554p 0 636.308p 0 636.309p 10000.0u 636.31p 0 637.415p 0 637.416p 10000.0u 637.417p 0 647.921p 0 647.922p 10000.0u 647.923p 0 656.945p 0 656.946p 10000.0u 656.947p 0 657.575p 0 657.576p 10000.0u 657.577p 0 669.566p 0 669.567p 10000.0u 669.568p 0 681.164p 0 681.165p 10000.0u 681.166p 0 688.988p 0 688.989p 10000.0u 688.99p 0 707.0p 0 707.001p 10000.0u 707.002p 0 721.199p 0 721.2p 10000.0u 721.201p 0 733.625p 0 733.626p 10000.0u 733.627p 0 734.189p 0 734.19p 10000.0u 734.191p 0 737.507p 0 737.508p 10000.0u 737.509p 0 740.213p 0 740.214p 10000.0u 740.215p 0 742.16p 0 742.161p 10000.0u 742.162p 0 754.589p 0 754.59p 10000.0u 754.591p 0 756.746p 0 756.747p 10000.0u 756.748p 0 780.398p 0 780.399p 10000.0u 780.4p 0 806.081p 0 806.082p 10000.0u 806.083p 0 806.867p 0 806.868p 10000.0u 806.869p 0 811.466p 0 811.467p 10000.0u 811.468p 0 839.618p 0 839.619p 10000.0u 839.62p 0 840.365p 0 840.366p 10000.0u 840.367p 0 846.368p 0 846.369p 10000.0u 846.37p 0 861.62p 0 861.621p 10000.0u 861.622p 0 867.734p 0 867.735p 10000.0u 867.736p 0 873.764p 0 873.765p 10000.0u 873.766p 0 895.982p 0 895.983p 10000.0u 895.984p 0 897.041p 0 897.042p 10000.0u 897.043p 0 904.991p 0 904.992p 10000.0u 904.993p 0 908.612p 0 908.613p 10000.0u 908.614p 0 922.499p 0 922.5p 10000.0u 922.501p 0 925.598p 0 925.599p 10000.0u 925.6p 0 926.213p 0 926.214p 10000.0u 926.215p 0 944.96p 0 944.961p 10000.0u 944.962p 0 951.485p 0 951.486p 10000.0u 951.487p 0 955.295p 0 955.296p 10000.0u 955.297p 0 957.383p 0 957.384p 10000.0u 957.385p 0 973.559p 0 973.56p 10000.0u 973.561p 0 975.623p 0 975.624p 10000.0u 975.625p 0 988.265p 0 988.266p 10000.0u 988.267p 0)
IIN28 0 29 pwl(0 0 18.491p 0 18.492p 10000.0u 18.493p 0 23.873p 0 23.874p 10000.0u 23.875p 0 32.399p 0 32.4p 10000.0u 32.401p 0 36.863p 0 36.864p 10000.0u 36.865p 0 41.063p 0 41.064p 10000.0u 41.065p 0 42.53p 0 42.531p 10000.0u 42.532p 0 81.92p 0 81.921p 10000.0u 81.922p 0 98.132p 0 98.133p 10000.0u 98.134p 0 111.482p 0 111.483p 10000.0u 111.484p 0 120.509p 0 120.51p 10000.0u 120.511p 0 133.223p 0 133.224p 10000.0u 133.225p 0 157.133p 0 157.134p 10000.0u 157.135p 0 169.715p 0 169.716p 10000.0u 169.717p 0 181.835p 0 181.836p 10000.0u 181.837p 0 183.227p 0 183.228p 10000.0u 183.229p 0 193.856p 0 193.857p 10000.0u 193.858p 0 195.17p 0 195.171p 10000.0u 195.172p 0 200.807p 0 200.808p 10000.0u 200.809p 0 246.989p 0 246.99p 10000.0u 246.991p 0 248.396p 0 248.397p 10000.0u 248.398p 0 252.509p 0 252.51p 10000.0u 252.511p 0 259.427p 0 259.428p 10000.0u 259.429p 0 267.083p 0 267.084p 10000.0u 267.085p 0 269.942p 0 269.943p 10000.0u 269.944p 0 269.972p 0 269.973p 10000.0u 269.974p 0 278.315p 0 278.316p 10000.0u 278.317p 0 285.5p 0 285.501p 10000.0u 285.502p 0 291.233p 0 291.234p 10000.0u 291.235p 0 302.501p 0 302.502p 10000.0u 302.503p 0 313.355p 0 313.356p 10000.0u 313.357p 0 348.707p 0 348.708p 10000.0u 348.709p 0 350.624p 0 350.625p 10000.0u 350.626p 0 373.328p 0 373.329p 10000.0u 373.33p 0 381.974p 0 381.975p 10000.0u 381.976p 0 388.076p 0 388.077p 10000.0u 388.078p 0 392.423p 0 392.424p 10000.0u 392.425p 0 398.723p 0 398.724p 10000.0u 398.725p 0 406.19p 0 406.191p 10000.0u 406.192p 0 416.72p 0 416.721p 10000.0u 416.722p 0 417.665p 0 417.666p 10000.0u 417.667p 0 421.601p 0 421.602p 10000.0u 421.603p 0 459.617p 0 459.618p 10000.0u 459.619p 0 465.071p 0 465.072p 10000.0u 465.073p 0 489.647p 0 489.648p 10000.0u 489.649p 0 494.348p 0 494.349p 10000.0u 494.35p 0 505.856p 0 505.857p 10000.0u 505.858p 0 506.756p 0 506.757p 10000.0u 506.758p 0 513.95p 0 513.951p 10000.0u 513.952p 0 518.753p 0 518.754p 10000.0u 518.755p 0 527.717p 0 527.718p 10000.0u 527.719p 0 528.581p 0 528.582p 10000.0u 528.583p 0 545.282p 0 545.283p 10000.0u 545.284p 0 567.131p 0 567.132p 10000.0u 567.133p 0 572.495p 0 572.496p 10000.0u 572.497p 0 573.53p 0 573.531p 10000.0u 573.532p 0 579.599p 0 579.6p 10000.0u 579.601p 0 585.605p 0 585.606p 10000.0u 585.607p 0 586.904p 0 586.905p 10000.0u 586.906p 0 607.475p 0 607.476p 10000.0u 607.477p 0 632.057p 0 632.058p 10000.0u 632.059p 0 641.633p 0 641.634p 10000.0u 641.635p 0 652.841p 0 652.842p 10000.0u 652.843p 0 658.814p 0 658.815p 10000.0u 658.816p 0 660.41p 0 660.411p 10000.0u 660.412p 0 665.447p 0 665.448p 10000.0u 665.449p 0 673.562p 0 673.563p 10000.0u 673.564p 0 681.71p 0 681.711p 10000.0u 681.712p 0 688.943p 0 688.944p 10000.0u 688.945p 0 705.779p 0 705.78p 10000.0u 705.781p 0 708.626p 0 708.627p 10000.0u 708.628p 0 732.509p 0 732.51p 10000.0u 732.511p 0 733.394p 0 733.395p 10000.0u 733.396p 0 737.042p 0 737.043p 10000.0u 737.044p 0 739.199p 0 739.2p 10000.0u 739.201p 0 742.433p 0 742.434p 10000.0u 742.435p 0 771.857p 0 771.858p 10000.0u 771.859p 0 776.348p 0 776.349p 10000.0u 776.35p 0 776.498p 0 776.499p 10000.0u 776.5p 0 785.945p 0 785.946p 10000.0u 785.947p 0 796.406p 0 796.407p 10000.0u 796.408p 0 800.591p 0 800.592p 10000.0u 800.593p 0 802.118p 0 802.119p 10000.0u 802.12p 0 806.372p 0 806.373p 10000.0u 806.374p 0 813.134p 0 813.135p 10000.0u 813.136p 0 819.716p 0 819.717p 10000.0u 819.718p 0 832.673p 0 832.674p 10000.0u 832.675p 0 840.488p 0 840.489p 10000.0u 840.49p 0 847.589p 0 847.59p 10000.0u 847.591p 0 900.023p 0 900.024p 10000.0u 900.025p 0 907.175p 0 907.176p 10000.0u 907.177p 0 911.51p 0 911.511p 10000.0u 911.512p 0 930.068p 0 930.069p 10000.0u 930.07p 0 941.498p 0 941.499p 10000.0u 941.5p 0 955.439p 0 955.44p 10000.0u 955.441p 0 962.876p 0 962.877p 10000.0u 962.878p 0 975.74p 0 975.741p 10000.0u 975.742p 0 995.597p 0 995.598p 10000.0u 995.599p 0 999.062p 0 999.063p 10000.0u 999.064p 0 999.434p 0 999.435p 10000.0u 999.436p 0)
IIN29 0 30 pwl(0 0 7.859p 0 7.86p 10000.0u 7.861p 0 25.508p 0 25.509p 10000.0u 25.51p 0 52.838p 0 52.839p 10000.0u 52.84p 0 59.825p 0 59.826p 10000.0u 59.827p 0 59.978p 0 59.979p 10000.0u 59.98p 0 61.136p 0 61.137p 10000.0u 61.138p 0 63.806p 0 63.807p 10000.0u 63.808p 0 89.135p 0 89.136p 10000.0u 89.137p 0 95.582p 0 95.583p 10000.0u 95.584p 0 100.325p 0 100.326p 10000.0u 100.327p 0 121.031p 0 121.032p 10000.0u 121.033p 0 132.011p 0 132.012p 10000.0u 132.013p 0 160.025p 0 160.026p 10000.0u 160.027p 0 173.258p 0 173.259p 10000.0u 173.26p 0 200.432p 0 200.433p 10000.0u 200.434p 0 218.213p 0 218.214p 10000.0u 218.215p 0 247.184p 0 247.185p 10000.0u 247.186p 0 250.961p 0 250.962p 10000.0u 250.963p 0 257.603p 0 257.604p 10000.0u 257.605p 0 259.619p 0 259.62p 10000.0u 259.621p 0 260.345p 0 260.346p 10000.0u 260.347p 0 278.783p 0 278.784p 10000.0u 278.785p 0 279.035p 0 279.036p 10000.0u 279.037p 0 281.903p 0 281.904p 10000.0u 281.905p 0 284.264p 0 284.265p 10000.0u 284.266p 0 284.741p 0 284.742p 10000.0u 284.743p 0 285.845p 0 285.846p 10000.0u 285.847p 0 291.197p 0 291.198p 10000.0u 291.199p 0 301.358p 0 301.359p 10000.0u 301.36p 0 312.617p 0 312.618p 10000.0u 312.619p 0 318.656p 0 318.657p 10000.0u 318.658p 0 319.457p 0 319.458p 10000.0u 319.459p 0 346.67p 0 346.671p 10000.0u 346.672p 0 348.554p 0 348.555p 10000.0u 348.556p 0 357.095p 0 357.096p 10000.0u 357.097p 0 371.564p 0 371.565p 10000.0u 371.566p 0 376.568p 0 376.569p 10000.0u 376.57p 0 382.835p 0 382.836p 10000.0u 382.837p 0 384.461p 0 384.462p 10000.0u 384.463p 0 384.695p 0 384.696p 10000.0u 384.697p 0 406.292p 0 406.293p 10000.0u 406.294p 0 459.008p 0 459.009p 10000.0u 459.01p 0 464.195p 0 464.196p 10000.0u 464.197p 0 464.204p 0 464.205p 10000.0u 464.206p 0 477.164p 0 477.165p 10000.0u 477.166p 0 488.582p 0 488.583p 10000.0u 488.584p 0 494.837p 0 494.838p 10000.0u 494.839p 0 518.864p 0 518.865p 10000.0u 518.866p 0 519.47p 0 519.471p 10000.0u 519.472p 0 524.84p 0 524.841p 10000.0u 524.842p 0 528.71p 0 528.711p 10000.0u 528.712p 0 528.956p 0 528.957p 10000.0u 528.958p 0 536.303p 0 536.304p 10000.0u 536.305p 0 544.265p 0 544.266p 10000.0u 544.267p 0 548.069p 0 548.07p 10000.0u 548.071p 0 560.294p 0 560.295p 10000.0u 560.296p 0 561.497p 0 561.498p 10000.0u 561.499p 0 604.079p 0 604.08p 10000.0u 604.081p 0 605.471p 0 605.472p 10000.0u 605.473p 0 609.038p 0 609.039p 10000.0u 609.04p 0 612.029p 0 612.03p 10000.0u 612.031p 0 616.145p 0 616.146p 10000.0u 616.147p 0 632.267p 0 632.268p 10000.0u 632.269p 0 650.252p 0 650.253p 10000.0u 650.254p 0 650.546p 0 650.547p 10000.0u 650.548p 0 655.247p 0 655.248p 10000.0u 655.249p 0 663.917p 0 663.918p 10000.0u 663.919p 0 665.102p 0 665.103p 10000.0u 665.104p 0 703.652p 0 703.653p 10000.0u 703.654p 0 716.096p 0 716.097p 10000.0u 716.098p 0 746.237p 0 746.238p 10000.0u 746.239p 0 752.615p 0 752.616p 10000.0u 752.617p 0 766.097p 0 766.098p 10000.0u 766.099p 0 766.496p 0 766.497p 10000.0u 766.498p 0 770.519p 0 770.52p 10000.0u 770.521p 0 776.108p 0 776.109p 10000.0u 776.11p 0 784.268p 0 784.269p 10000.0u 784.27p 0 786.743p 0 786.744p 10000.0u 786.745p 0 793.691p 0 793.692p 10000.0u 793.693p 0 801.674p 0 801.675p 10000.0u 801.676p 0 806.507p 0 806.508p 10000.0u 806.509p 0 814.958p 0 814.959p 10000.0u 814.96p 0 823.013p 0 823.014p 10000.0u 823.015p 0 830.711p 0 830.712p 10000.0u 830.713p 0 835.355p 0 835.356p 10000.0u 835.357p 0 848.969p 0 848.97p 10000.0u 848.971p 0 851.492p 0 851.493p 10000.0u 851.494p 0 862.829p 0 862.83p 10000.0u 862.831p 0 874.856p 0 874.857p 10000.0u 874.858p 0 880.622p 0 880.623p 10000.0u 880.624p 0 881.288p 0 881.289p 10000.0u 881.29p 0 881.717p 0 881.718p 10000.0u 881.719p 0 885.827p 0 885.828p 10000.0u 885.829p 0 901.697p 0 901.698p 10000.0u 901.699p 0 911.741p 0 911.742p 10000.0u 911.743p 0 923.327p 0 923.328p 10000.0u 923.329p 0 931.166p 0 931.167p 10000.0u 931.168p 0 966.173p 0 966.174p 10000.0u 966.175p 0 966.599p 0 966.6p 10000.0u 966.601p 0 966.986p 0 966.987p 10000.0u 966.988p 0 972.35p 0 972.351p 10000.0u 972.352p 0)
IIN30 0 31 pwl(0 0 4.388p 0 4.389p 10000.0u 4.39p 0 18.551p 0 18.552p 10000.0u 18.553p 0 24.338p 0 24.339p 10000.0u 24.34p 0 36.467p 0 36.468p 10000.0u 36.469p 0 79.223p 0 79.224p 10000.0u 79.225p 0 81.824p 0 81.825p 10000.0u 81.826p 0 113.819p 0 113.82p 10000.0u 113.821p 0 117.644p 0 117.645p 10000.0u 117.646p 0 122.639p 0 122.64p 10000.0u 122.641p 0 138.011p 0 138.012p 10000.0u 138.013p 0 176.792p 0 176.793p 10000.0u 176.794p 0 202.307p 0 202.308p 10000.0u 202.309p 0 207.266p 0 207.267p 10000.0u 207.268p 0 223.961p 0 223.962p 10000.0u 223.963p 0 227.861p 0 227.862p 10000.0u 227.863p 0 231.059p 0 231.06p 10000.0u 231.061p 0 233.66p 0 233.661p 10000.0u 233.662p 0 236.408p 0 236.409p 10000.0u 236.41p 0 238.667p 0 238.668p 10000.0u 238.669p 0 292.289p 0 292.29p 10000.0u 292.291p 0 304.154p 0 304.155p 10000.0u 304.156p 0 326.264p 0 326.265p 10000.0u 326.266p 0 327.335p 0 327.336p 10000.0u 327.337p 0 335.369p 0 335.37p 10000.0u 335.371p 0 344.537p 0 344.538p 10000.0u 344.539p 0 351.641p 0 351.642p 10000.0u 351.643p 0 352.31p 0 352.311p 10000.0u 352.312p 0 375.284p 0 375.285p 10000.0u 375.286p 0 395.684p 0 395.685p 10000.0u 395.686p 0 400.913p 0 400.914p 10000.0u 400.915p 0 430.601p 0 430.602p 10000.0u 430.603p 0 441.188p 0 441.189p 10000.0u 441.19p 0 448.448p 0 448.449p 10000.0u 448.45p 0 448.463p 0 448.464p 10000.0u 448.465p 0 448.901p 0 448.902p 10000.0u 448.903p 0 449.069p 0 449.07p 10000.0u 449.071p 0 452.525p 0 452.526p 10000.0u 452.527p 0 460.139p 0 460.14p 10000.0u 460.141p 0 474.053p 0 474.054p 10000.0u 474.055p 0 474.908p 0 474.909p 10000.0u 474.91p 0 494.12p 0 494.121p 10000.0u 494.122p 0 518.963p 0 518.964p 10000.0u 518.965p 0 519.431p 0 519.432p 10000.0u 519.433p 0 519.842p 0 519.843p 10000.0u 519.844p 0 525.314p 0 525.315p 10000.0u 525.316p 0 526.091p 0 526.092p 10000.0u 526.093p 0 550.7p 0 550.701p 10000.0u 550.702p 0 554.771p 0 554.772p 10000.0u 554.773p 0 556.475p 0 556.476p 10000.0u 556.477p 0 567.881p 0 567.882p 10000.0u 567.883p 0 568.505p 0 568.506p 10000.0u 568.507p 0 588.578p 0 588.579p 10000.0u 588.58p 0 591.71p 0 591.711p 10000.0u 591.712p 0 593.42p 0 593.421p 10000.0u 593.422p 0 613.322p 0 613.323p 10000.0u 613.324p 0 618.794p 0 618.795p 10000.0u 618.796p 0 622.199p 0 622.2p 10000.0u 622.201p 0 627.665p 0 627.666p 10000.0u 627.667p 0 629.03p 0 629.031p 10000.0u 629.032p 0 638.759p 0 638.76p 10000.0u 638.761p 0 639.734p 0 639.735p 10000.0u 639.736p 0 640.178p 0 640.179p 10000.0u 640.18p 0 641.864p 0 641.865p 10000.0u 641.866p 0 654.674p 0 654.675p 10000.0u 654.676p 0 660.146p 0 660.147p 10000.0u 660.148p 0 665.537p 0 665.538p 10000.0u 665.539p 0 673.145p 0 673.146p 10000.0u 673.147p 0 689.357p 0 689.358p 10000.0u 689.359p 0 695.231p 0 695.232p 10000.0u 695.233p 0 704.027p 0 704.028p 10000.0u 704.029p 0 711.353p 0 711.354p 10000.0u 711.355p 0 711.854p 0 711.855p 10000.0u 711.856p 0 720.116p 0 720.117p 10000.0u 720.118p 0 723.821p 0 723.822p 10000.0u 723.823p 0 729.638p 0 729.639p 10000.0u 729.64p 0 744.527p 0 744.528p 10000.0u 744.529p 0 761.882p 0 761.883p 10000.0u 761.884p 0 763.415p 0 763.416p 10000.0u 763.417p 0 767.03p 0 767.031p 10000.0u 767.032p 0 779.45p 0 779.451p 10000.0u 779.452p 0 793.733p 0 793.734p 10000.0u 793.735p 0 826.838p 0 826.839p 10000.0u 826.84p 0 828.722p 0 828.723p 10000.0u 828.724p 0 830.084p 0 830.085p 10000.0u 830.086p 0 861.344p 0 861.345p 10000.0u 861.346p 0 862.592p 0 862.593p 10000.0u 862.594p 0 886.34p 0 886.341p 10000.0u 886.342p 0 896.579p 0 896.58p 10000.0u 896.581p 0 898.544p 0 898.545p 10000.0u 898.546p 0 903.236p 0 903.237p 10000.0u 903.238p 0 905.417p 0 905.418p 10000.0u 905.419p 0 911.069p 0 911.07p 10000.0u 911.071p 0 936.326p 0 936.327p 10000.0u 936.328p 0 937.364p 0 937.365p 10000.0u 937.366p 0 944.06p 0 944.061p 10000.0u 944.062p 0 953.399p 0 953.4p 10000.0u 953.401p 0 965.474p 0 965.475p 10000.0u 965.476p 0 973.619p 0 973.62p 10000.0u 973.621p 0 973.688p 0 973.689p 10000.0u 973.69p 0 976.181p 0 976.182p 10000.0u 976.183p 0 977.63p 0 977.631p 10000.0u 977.632p 0 977.903p 0 977.904p 10000.0u 977.905p 0 979.847p 0 979.848p 10000.0u 979.849p 0 981.536p 0 981.537p 10000.0u 981.538p 0 986.027p 0 986.028p 10000.0u 986.029p 0 988.823p 0 988.824p 10000.0u 988.825p 0 995.39p 0 995.391p 10000.0u 995.392p 0)
IIN31 0 32 pwl(0 0 34.052p 0 34.053p 10000.0u 34.054p 0 36.359p 0 36.36p 10000.0u 36.361p 0 36.767p 0 36.768p 10000.0u 36.769p 0 41.321p 0 41.322p 10000.0u 41.323p 0 43.745p 0 43.746p 10000.0u 43.747p 0 52.277p 0 52.278p 10000.0u 52.279p 0 54.128p 0 54.129p 10000.0u 54.13p 0 58.187p 0 58.188p 10000.0u 58.189p 0 69.293p 0 69.294p 10000.0u 69.295p 0 81.035p 0 81.036p 10000.0u 81.037p 0 82.328p 0 82.329p 10000.0u 82.33p 0 94.424p 0 94.425p 10000.0u 94.426p 0 96.506p 0 96.507p 10000.0u 96.508p 0 118.031p 0 118.032p 10000.0u 118.033p 0 118.172p 0 118.173p 10000.0u 118.174p 0 125.897p 0 125.898p 10000.0u 125.899p 0 136.907p 0 136.908p 10000.0u 136.909p 0 139.046p 0 139.047p 10000.0u 139.048p 0 139.262p 0 139.263p 10000.0u 139.264p 0 144.47p 0 144.471p 10000.0u 144.472p 0 162.734p 0 162.735p 10000.0u 162.736p 0 172.595p 0 172.596p 10000.0u 172.597p 0 174.119p 0 174.12p 10000.0u 174.121p 0 174.863p 0 174.864p 10000.0u 174.865p 0 177.413p 0 177.414p 10000.0u 177.415p 0 189.194p 0 189.195p 10000.0u 189.196p 0 190.901p 0 190.902p 10000.0u 190.903p 0 197.15p 0 197.151p 10000.0u 197.152p 0 201.194p 0 201.195p 10000.0u 201.196p 0 205.343p 0 205.344p 10000.0u 205.345p 0 218.663p 0 218.664p 10000.0u 218.665p 0 224.885p 0 224.886p 10000.0u 224.887p 0 225.803p 0 225.804p 10000.0u 225.805p 0 243.158p 0 243.159p 10000.0u 243.16p 0 257.945p 0 257.946p 10000.0u 257.947p 0 269.111p 0 269.112p 10000.0u 269.113p 0 269.597p 0 269.598p 10000.0u 269.599p 0 276.851p 0 276.852p 10000.0u 276.853p 0 281.261p 0 281.262p 10000.0u 281.263p 0 285.557p 0 285.558p 10000.0u 285.559p 0 298.859p 0 298.86p 10000.0u 298.861p 0 304.049p 0 304.05p 10000.0u 304.051p 0 333.896p 0 333.897p 10000.0u 333.898p 0 342.914p 0 342.915p 10000.0u 342.916p 0 367.793p 0 367.794p 10000.0u 367.795p 0 379.034p 0 379.035p 10000.0u 379.036p 0 393.146p 0 393.147p 10000.0u 393.148p 0 395.03p 0 395.031p 10000.0u 395.032p 0 432.629p 0 432.63p 10000.0u 432.631p 0 453.872p 0 453.873p 10000.0u 453.874p 0 454.814p 0 454.815p 10000.0u 454.816p 0 484.694p 0 484.695p 10000.0u 484.696p 0 490.844p 0 490.845p 10000.0u 490.846p 0 509.549p 0 509.55p 10000.0u 509.551p 0 512.672p 0 512.673p 10000.0u 512.674p 0 514.271p 0 514.272p 10000.0u 514.273p 0 525.599p 0 525.6p 10000.0u 525.601p 0 532.082p 0 532.083p 10000.0u 532.084p 0 554.681p 0 554.682p 10000.0u 554.683p 0 557.936p 0 557.937p 10000.0u 557.938p 0 586.907p 0 586.908p 10000.0u 586.909p 0 588.293p 0 588.294p 10000.0u 588.295p 0 608.294p 0 608.295p 10000.0u 608.296p 0 640.61p 0 640.611p 10000.0u 640.612p 0 659.141p 0 659.142p 10000.0u 659.143p 0 668.417p 0 668.418p 10000.0u 668.419p 0 678.428p 0 678.429p 10000.0u 678.43p 0 681.488p 0 681.489p 10000.0u 681.49p 0 691.739p 0 691.74p 10000.0u 691.741p 0 708.809p 0 708.81p 10000.0u 708.811p 0 710.729p 0 710.73p 10000.0u 710.731p 0 724.148p 0 724.149p 10000.0u 724.15p 0 726.593p 0 726.594p 10000.0u 726.595p 0 727.577p 0 727.578p 10000.0u 727.579p 0 732.575p 0 732.576p 10000.0u 732.577p 0 743.888p 0 743.889p 10000.0u 743.89p 0 749.645p 0 749.646p 10000.0u 749.647p 0 751.568p 0 751.569p 10000.0u 751.57p 0 776.777p 0 776.778p 10000.0u 776.779p 0 777.572p 0 777.573p 10000.0u 777.574p 0 788.501p 0 788.502p 10000.0u 788.503p 0 799.445p 0 799.446p 10000.0u 799.447p 0 809.426p 0 809.427p 10000.0u 809.428p 0 828.008p 0 828.009p 10000.0u 828.01p 0 836.825p 0 836.826p 10000.0u 836.827p 0 860.294p 0 860.295p 10000.0u 860.296p 0 865.52p 0 865.521p 10000.0u 865.522p 0 866.666p 0 866.667p 10000.0u 866.668p 0 870.881p 0 870.882p 10000.0u 870.883p 0 889.742p 0 889.743p 10000.0u 889.744p 0 895.361p 0 895.362p 10000.0u 895.363p 0 943.394p 0 943.395p 10000.0u 943.396p 0 947.579p 0 947.58p 10000.0u 947.581p 0 959.081p 0 959.082p 10000.0u 959.083p 0 971.144p 0 971.145p 10000.0u 971.146p 0 992.738p 0 992.739p 10000.0u 992.74p 0 997.826p 0 997.827p 10000.0u 997.828p 0)
IIN32 0 33 pwl(0 0 13.367p 0 13.368p 10000.0u 13.369p 0 13.682p 0 13.683p 10000.0u 13.684p 0 16.073p 0 16.074p 10000.0u 16.075p 0 22.799p 0 22.8p 10000.0u 22.801p 0 27.044p 0 27.045p 10000.0u 27.046p 0 41.228p 0 41.229p 10000.0u 41.23p 0 51.974p 0 51.975p 10000.0u 51.976p 0 55.364p 0 55.365p 10000.0u 55.366p 0 59.414p 0 59.415p 10000.0u 59.416p 0 60.329p 0 60.33p 10000.0u 60.331p 0 60.875p 0 60.876p 10000.0u 60.877p 0 85.064p 0 85.065p 10000.0u 85.066p 0 89.357p 0 89.358p 10000.0u 89.359p 0 90.143p 0 90.144p 10000.0u 90.145p 0 132.44p 0 132.441p 10000.0u 132.442p 0 136.592p 0 136.593p 10000.0u 136.594p 0 139.421p 0 139.422p 10000.0u 139.423p 0 150.575p 0 150.576p 10000.0u 150.577p 0 169.211p 0 169.212p 10000.0u 169.213p 0 174.431p 0 174.432p 10000.0u 174.433p 0 184.835p 0 184.836p 10000.0u 184.837p 0 223.517p 0 223.518p 10000.0u 223.519p 0 237.212p 0 237.213p 10000.0u 237.214p 0 239.096p 0 239.097p 10000.0u 239.098p 0 244.328p 0 244.329p 10000.0u 244.33p 0 252.464p 0 252.465p 10000.0u 252.466p 0 254.225p 0 254.226p 10000.0u 254.227p 0 260.939p 0 260.94p 10000.0u 260.941p 0 267.992p 0 267.993p 10000.0u 267.994p 0 285.77p 0 285.771p 10000.0u 285.772p 0 294.713p 0 294.714p 10000.0u 294.715p 0 315.458p 0 315.459p 10000.0u 315.46p 0 319.871p 0 319.872p 10000.0u 319.873p 0 324.569p 0 324.57p 10000.0u 324.571p 0 327.848p 0 327.849p 10000.0u 327.85p 0 328.01p 0 328.011p 10000.0u 328.012p 0 334.289p 0 334.29p 10000.0u 334.291p 0 334.7p 0 334.701p 10000.0u 334.702p 0 345.446p 0 345.447p 10000.0u 345.448p 0 350.237p 0 350.238p 10000.0u 350.239p 0 352.319p 0 352.32p 10000.0u 352.321p 0 355.046p 0 355.047p 10000.0u 355.048p 0 390.446p 0 390.447p 10000.0u 390.448p 0 401.6p 0 401.601p 10000.0u 401.602p 0 415.145p 0 415.146p 10000.0u 415.147p 0 416.249p 0 416.25p 10000.0u 416.251p 0 451.298p 0 451.299p 10000.0u 451.3p 0 454.313p 0 454.314p 10000.0u 454.315p 0 467.219p 0 467.22p 10000.0u 467.221p 0 467.783p 0 467.784p 10000.0u 467.785p 0 470.657p 0 470.658p 10000.0u 470.659p 0 476.537p 0 476.538p 10000.0u 476.539p 0 478.037p 0 478.038p 10000.0u 478.039p 0 485.009p 0 485.01p 10000.0u 485.011p 0 546.323p 0 546.324p 10000.0u 546.325p 0 555.614p 0 555.615p 10000.0u 555.616p 0 633.587p 0 633.588p 10000.0u 633.589p 0 640.295p 0 640.296p 10000.0u 640.297p 0 645.476p 0 645.477p 10000.0u 645.478p 0 645.551p 0 645.552p 10000.0u 645.553p 0 650.705p 0 650.706p 10000.0u 650.707p 0 650.768p 0 650.769p 10000.0u 650.77p 0 664.7p 0 664.701p 10000.0u 664.702p 0 670.007p 0 670.008p 10000.0u 670.009p 0 671.774p 0 671.775p 10000.0u 671.776p 0 674.0p 0 674.001p 10000.0u 674.002p 0 678.89p 0 678.891p 10000.0u 678.892p 0 679.292p 0 679.293p 10000.0u 679.294p 0 696.209p 0 696.21p 10000.0u 696.211p 0 696.626p 0 696.627p 10000.0u 696.628p 0 709.541p 0 709.542p 10000.0u 709.543p 0 715.037p 0 715.038p 10000.0u 715.039p 0 718.616p 0 718.617p 10000.0u 718.618p 0 719.621p 0 719.622p 10000.0u 719.623p 0 720.221p 0 720.222p 10000.0u 720.223p 0 733.097p 0 733.098p 10000.0u 733.099p 0 764.327p 0 764.328p 10000.0u 764.329p 0 765.254p 0 765.255p 10000.0u 765.256p 0 769.088p 0 769.089p 10000.0u 769.09p 0 783.497p 0 783.498p 10000.0u 783.499p 0 811.058p 0 811.059p 10000.0u 811.06p 0 835.841p 0 835.842p 10000.0u 835.843p 0 837.389p 0 837.39p 10000.0u 837.391p 0 845.699p 0 845.7p 10000.0u 845.701p 0 865.994p 0 865.995p 10000.0u 865.996p 0 873.584p 0 873.585p 10000.0u 873.586p 0 892.871p 0 892.872p 10000.0u 892.873p 0 898.427p 0 898.428p 10000.0u 898.429p 0 916.394p 0 916.395p 10000.0u 916.396p 0 918.104p 0 918.105p 10000.0u 918.106p 0 920.828p 0 920.829p 10000.0u 920.83p 0 933.371p 0 933.372p 10000.0u 933.373p 0 936.833p 0 936.834p 10000.0u 936.835p 0 937.076p 0 937.077p 10000.0u 937.078p 0 943.856p 0 943.857p 10000.0u 943.858p 0 945.188p 0 945.189p 10000.0u 945.19p 0 954.848p 0 954.849p 10000.0u 954.85p 0 958.256p 0 958.257p 10000.0u 958.258p 0 976.181p 0 976.182p 10000.0u 976.183p 0 983.312p 0 983.313p 10000.0u 983.314p 0)
IIN33 0 34 pwl(0 0 1.646p 0 1.647p 10000.0u 1.648p 0 24.14p 0 24.141p 10000.0u 24.142p 0 25.475p 0 25.476p 10000.0u 25.477p 0 53.201p 0 53.202p 10000.0u 53.203p 0 54.881p 0 54.882p 10000.0u 54.883p 0 79.61p 0 79.611p 10000.0u 79.612p 0 89.48p 0 89.481p 10000.0u 89.482p 0 89.921p 0 89.922p 10000.0u 89.923p 0 93.383p 0 93.384p 10000.0u 93.385p 0 97.457p 0 97.458p 10000.0u 97.459p 0 102.566p 0 102.567p 10000.0u 102.568p 0 108.254p 0 108.255p 10000.0u 108.256p 0 122.396p 0 122.397p 10000.0u 122.398p 0 132.02p 0 132.021p 10000.0u 132.022p 0 133.301p 0 133.302p 10000.0u 133.303p 0 136.19p 0 136.191p 10000.0u 136.192p 0 141.752p 0 141.753p 10000.0u 141.754p 0 145.181p 0 145.182p 10000.0u 145.183p 0 147.896p 0 147.897p 10000.0u 147.898p 0 151.889p 0 151.89p 10000.0u 151.891p 0 182.414p 0 182.415p 10000.0u 182.416p 0 189.509p 0 189.51p 10000.0u 189.511p 0 190.139p 0 190.14p 10000.0u 190.141p 0 202.241p 0 202.242p 10000.0u 202.243p 0 203.606p 0 203.607p 10000.0u 203.608p 0 222.095p 0 222.096p 10000.0u 222.097p 0 227.705p 0 227.706p 10000.0u 227.707p 0 262.943p 0 262.944p 10000.0u 262.945p 0 269.438p 0 269.439p 10000.0u 269.44p 0 270.584p 0 270.585p 10000.0u 270.586p 0 274.499p 0 274.5p 10000.0u 274.501p 0 286.271p 0 286.272p 10000.0u 286.273p 0 287.693p 0 287.694p 10000.0u 287.695p 0 301.505p 0 301.506p 10000.0u 301.507p 0 310.181p 0 310.182p 10000.0u 310.183p 0 319.346p 0 319.347p 10000.0u 319.348p 0 328.145p 0 328.146p 10000.0u 328.147p 0 339.185p 0 339.186p 10000.0u 339.187p 0 349.466p 0 349.467p 10000.0u 349.468p 0 350.336p 0 350.337p 10000.0u 350.338p 0 361.328p 0 361.329p 10000.0u 361.33p 0 370.34p 0 370.341p 10000.0u 370.342p 0 380.393p 0 380.394p 10000.0u 380.395p 0 386.441p 0 386.442p 10000.0u 386.443p 0 416.441p 0 416.442p 10000.0u 416.443p 0 418.979p 0 418.98p 10000.0u 418.981p 0 423.332p 0 423.333p 10000.0u 423.334p 0 447.704p 0 447.705p 10000.0u 447.706p 0 450.008p 0 450.009p 10000.0u 450.01p 0 450.32p 0 450.321p 10000.0u 450.322p 0 454.538p 0 454.539p 10000.0u 454.54p 0 466.994p 0 466.995p 10000.0u 466.996p 0 481.151p 0 481.152p 10000.0u 481.153p 0 486.77p 0 486.771p 10000.0u 486.772p 0 495.968p 0 495.969p 10000.0u 495.97p 0 524.606p 0 524.607p 10000.0u 524.608p 0 526.322p 0 526.323p 10000.0u 526.324p 0 532.625p 0 532.626p 10000.0u 532.627p 0 549.752p 0 549.753p 10000.0u 549.754p 0 554.27p 0 554.271p 10000.0u 554.272p 0 557.585p 0 557.586p 10000.0u 557.587p 0 576.593p 0 576.594p 10000.0u 576.595p 0 576.758p 0 576.759p 10000.0u 576.76p 0 579.059p 0 579.06p 10000.0u 579.061p 0 584.174p 0 584.175p 10000.0u 584.176p 0 589.208p 0 589.209p 10000.0u 589.21p 0 590.807p 0 590.808p 10000.0u 590.809p 0 609.419p 0 609.42p 10000.0u 609.421p 0 620.552p 0 620.553p 10000.0u 620.554p 0 639.887p 0 639.888p 10000.0u 639.889p 0 659.057p 0 659.058p 10000.0u 659.059p 0 679.463p 0 679.464p 10000.0u 679.465p 0 692.843p 0 692.844p 10000.0u 692.845p 0 719.522p 0 719.523p 10000.0u 719.524p 0 720.377p 0 720.378p 10000.0u 720.379p 0 730.496p 0 730.497p 10000.0u 730.498p 0 732.821p 0 732.822p 10000.0u 732.823p 0 733.208p 0 733.209p 10000.0u 733.21p 0 738.53p 0 738.531p 10000.0u 738.532p 0 755.42p 0 755.421p 10000.0u 755.422p 0 756.38p 0 756.381p 10000.0u 756.382p 0 767.63p 0 767.631p 10000.0u 767.632p 0 774.344p 0 774.345p 10000.0u 774.346p 0 781.784p 0 781.785p 10000.0u 781.786p 0 785.492p 0 785.493p 10000.0u 785.494p 0 804.917p 0 804.918p 10000.0u 804.919p 0 820.58p 0 820.581p 10000.0u 820.582p 0 831.965p 0 831.966p 10000.0u 831.967p 0 832.649p 0 832.65p 10000.0u 832.651p 0 837.398p 0 837.399p 10000.0u 837.4p 0 868.907p 0 868.908p 10000.0u 868.909p 0 881.495p 0 881.496p 10000.0u 881.497p 0 883.826p 0 883.827p 10000.0u 883.828p 0 889.721p 0 889.722p 10000.0u 889.723p 0 891.248p 0 891.249p 10000.0u 891.25p 0 893.375p 0 893.376p 10000.0u 893.377p 0 911.519p 0 911.52p 10000.0u 911.521p 0 915.011p 0 915.012p 10000.0u 915.013p 0 919.139p 0 919.14p 10000.0u 919.141p 0 940.757p 0 940.758p 10000.0u 940.759p 0 942.536p 0 942.537p 10000.0u 942.538p 0 942.668p 0 942.669p 10000.0u 942.67p 0 965.252p 0 965.253p 10000.0u 965.254p 0 981.524p 0 981.525p 10000.0u 981.526p 0)
IIN34 0 35 pwl(0 0 6.218p 0 6.219p 10000.0u 6.22p 0 11.441p 0 11.442p 10000.0u 11.443p 0 20.828p 0 20.829p 10000.0u 20.83p 0 24.278p 0 24.279p 10000.0u 24.28p 0 44.588p 0 44.589p 10000.0u 44.59p 0 65.105p 0 65.106p 10000.0u 65.107p 0 90.785p 0 90.786p 10000.0u 90.787p 0 92.159p 0 92.16p 10000.0u 92.161p 0 108.554p 0 108.555p 10000.0u 108.556p 0 118.013p 0 118.014p 10000.0u 118.015p 0 137.873p 0 137.874p 10000.0u 137.875p 0 143.39p 0 143.391p 10000.0u 143.392p 0 175.604p 0 175.605p 10000.0u 175.606p 0 179.258p 0 179.259p 10000.0u 179.26p 0 189.332p 0 189.333p 10000.0u 189.334p 0 192.989p 0 192.99p 10000.0u 192.991p 0 203.432p 0 203.433p 10000.0u 203.434p 0 204.485p 0 204.486p 10000.0u 204.487p 0 210.386p 0 210.387p 10000.0u 210.388p 0 225.896p 0 225.897p 10000.0u 225.898p 0 230.573p 0 230.574p 10000.0u 230.575p 0 244.532p 0 244.533p 10000.0u 244.534p 0 250.445p 0 250.446p 10000.0u 250.447p 0 259.886p 0 259.887p 10000.0u 259.888p 0 267.755p 0 267.756p 10000.0u 267.757p 0 273.32p 0 273.321p 10000.0u 273.322p 0 277.058p 0 277.059p 10000.0u 277.06p 0 301.139p 0 301.14p 10000.0u 301.141p 0 332.282p 0 332.283p 10000.0u 332.284p 0 335.453p 0 335.454p 10000.0u 335.455p 0 338.048p 0 338.049p 10000.0u 338.05p 0 353.855p 0 353.856p 10000.0u 353.857p 0 355.655p 0 355.656p 10000.0u 355.657p 0 361.79p 0 361.791p 10000.0u 361.792p 0 371.627p 0 371.628p 10000.0u 371.629p 0 374.525p 0 374.526p 10000.0u 374.527p 0 389.066p 0 389.067p 10000.0u 389.068p 0 402.773p 0 402.774p 10000.0u 402.775p 0 410.933p 0 410.934p 10000.0u 410.935p 0 421.982p 0 421.983p 10000.0u 421.984p 0 452.729p 0 452.73p 10000.0u 452.731p 0 474.026p 0 474.027p 10000.0u 474.028p 0 479.411p 0 479.412p 10000.0u 479.413p 0 514.733p 0 514.734p 10000.0u 514.735p 0 520.781p 0 520.782p 10000.0u 520.783p 0 528.629p 0 528.63p 10000.0u 528.631p 0 539.876p 0 539.877p 10000.0u 539.878p 0 545.381p 0 545.382p 10000.0u 545.383p 0 555.269p 0 555.27p 10000.0u 555.271p 0 556.088p 0 556.089p 10000.0u 556.09p 0 558.479p 0 558.48p 10000.0u 558.481p 0 568.109p 0 568.11p 10000.0u 568.111p 0 575.195p 0 575.196p 10000.0u 575.197p 0 592.679p 0 592.68p 10000.0u 592.681p 0 602.75p 0 602.751p 10000.0u 602.752p 0 629.801p 0 629.802p 10000.0u 629.803p 0 635.12p 0 635.121p 10000.0u 635.122p 0 640.295p 0 640.296p 10000.0u 640.297p 0 645.659p 0 645.66p 10000.0u 645.661p 0 651.881p 0 651.882p 10000.0u 651.883p 0 653.363p 0 653.364p 10000.0u 653.365p 0 658.898p 0 658.899p 10000.0u 658.9p 0 661.115p 0 661.116p 10000.0u 661.117p 0 694.682p 0 694.683p 10000.0u 694.684p 0 727.946p 0 727.947p 10000.0u 727.948p 0 736.673p 0 736.674p 10000.0u 736.675p 0 736.94p 0 736.941p 10000.0u 736.942p 0 745.238p 0 745.239p 10000.0u 745.24p 0 753.533p 0 753.534p 10000.0u 753.535p 0 753.566p 0 753.567p 10000.0u 753.568p 0 755.891p 0 755.892p 10000.0u 755.893p 0 760.43p 0 760.431p 10000.0u 760.432p 0 790.076p 0 790.077p 10000.0u 790.078p 0 793.655p 0 793.656p 10000.0u 793.657p 0 793.724p 0 793.725p 10000.0u 793.726p 0 827.447p 0 827.448p 10000.0u 827.449p 0 828.551p 0 828.552p 10000.0u 828.553p 0 833.87p 0 833.871p 10000.0u 833.872p 0 839.981p 0 839.982p 10000.0u 839.983p 0 844.115p 0 844.116p 10000.0u 844.117p 0 845.261p 0 845.262p 10000.0u 845.263p 0 857.588p 0 857.589p 10000.0u 857.59p 0 870.014p 0 870.015p 10000.0u 870.016p 0 903.53p 0 903.531p 10000.0u 903.532p 0 910.28p 0 910.281p 10000.0u 910.282p 0 923.978p 0 923.979p 10000.0u 923.98p 0 926.111p 0 926.112p 10000.0u 926.113p 0 952.13p 0 952.131p 10000.0u 952.132p 0 955.055p 0 955.056p 10000.0u 955.057p 0 958.277p 0 958.278p 10000.0u 958.279p 0 983.921p 0 983.922p 10000.0u 983.923p 0 999.593p 0 999.594p 10000.0u 999.595p 0 999.677p 0 999.678p 10000.0u 999.679p 0)
IIN35 0 36 pwl(0 0 3.155p 0 3.156p 10000.0u 3.157p 0 5.264p 0 5.265p 10000.0u 5.266p 0 16.895p 0 16.896p 10000.0u 16.897p 0 17.096p 0 17.097p 10000.0u 17.098p 0 30.572p 0 30.573p 10000.0u 30.574p 0 33.575p 0 33.576p 10000.0u 33.577p 0 36.422p 0 36.423p 10000.0u 36.424p 0 45.926p 0 45.927p 10000.0u 45.928p 0 52.319p 0 52.32p 10000.0u 52.321p 0 59.807p 0 59.808p 10000.0u 59.809p 0 63.971p 0 63.972p 10000.0u 63.973p 0 74.351p 0 74.352p 10000.0u 74.353p 0 86.447p 0 86.448p 10000.0u 86.449p 0 88.529p 0 88.53p 10000.0u 88.531p 0 121.697p 0 121.698p 10000.0u 121.699p 0 124.757p 0 124.758p 10000.0u 124.759p 0 142.337p 0 142.338p 10000.0u 142.339p 0 142.472p 0 142.473p 10000.0u 142.474p 0 170.018p 0 170.019p 10000.0u 170.02p 0 184.808p 0 184.809p 10000.0u 184.81p 0 192.266p 0 192.267p 10000.0u 192.268p 0 198.995p 0 198.996p 10000.0u 198.997p 0 199.724p 0 199.725p 10000.0u 199.726p 0 205.226p 0 205.227p 10000.0u 205.228p 0 221.612p 0 221.613p 10000.0u 221.614p 0 237.299p 0 237.3p 10000.0u 237.301p 0 251.018p 0 251.019p 10000.0u 251.02p 0 264.977p 0 264.978p 10000.0u 264.979p 0 272.0p 0 272.001p 10000.0u 272.002p 0 272.972p 0 272.973p 10000.0u 272.974p 0 297.122p 0 297.123p 10000.0u 297.124p 0 315.314p 0 315.315p 10000.0u 315.316p 0 331.58p 0 331.581p 10000.0u 331.582p 0 334.874p 0 334.875p 10000.0u 334.876p 0 339.686p 0 339.687p 10000.0u 339.688p 0 351.413p 0 351.414p 10000.0u 351.415p 0 368.357p 0 368.358p 10000.0u 368.359p 0 374.108p 0 374.109p 10000.0u 374.11p 0 377.459p 0 377.46p 10000.0u 377.461p 0 397.127p 0 397.128p 10000.0u 397.129p 0 401.39p 0 401.391p 10000.0u 401.392p 0 401.681p 0 401.682p 10000.0u 401.683p 0 406.694p 0 406.695p 10000.0u 406.696p 0 449.627p 0 449.628p 10000.0u 449.629p 0 456.431p 0 456.432p 10000.0u 456.433p 0 461.552p 0 461.553p 10000.0u 461.554p 0 475.571p 0 475.572p 10000.0u 475.573p 0 475.757p 0 475.758p 10000.0u 475.759p 0 482.357p 0 482.358p 10000.0u 482.359p 0 503.201p 0 503.202p 10000.0u 503.203p 0 504.557p 0 504.558p 10000.0u 504.559p 0 509.768p 0 509.769p 10000.0u 509.77p 0 511.271p 0 511.272p 10000.0u 511.273p 0 520.895p 0 520.896p 10000.0u 520.897p 0 526.919p 0 526.92p 10000.0u 526.921p 0 538.238p 0 538.239p 10000.0u 538.24p 0 542.795p 0 542.796p 10000.0u 542.797p 0 546.968p 0 546.969p 10000.0u 546.97p 0 552.242p 0 552.243p 10000.0u 552.244p 0 554.444p 0 554.445p 10000.0u 554.446p 0 554.888p 0 554.889p 10000.0u 554.89p 0 564.359p 0 564.36p 10000.0u 564.361p 0 568.238p 0 568.239p 10000.0u 568.24p 0 569.195p 0 569.196p 10000.0u 569.197p 0 580.01p 0 580.011p 10000.0u 580.012p 0 614.537p 0 614.538p 10000.0u 614.539p 0 620.108p 0 620.109p 10000.0u 620.11p 0 625.433p 0 625.434p 10000.0u 625.435p 0 628.013p 0 628.014p 10000.0u 628.015p 0 628.601p 0 628.602p 10000.0u 628.603p 0 630.725p 0 630.726p 10000.0u 630.727p 0 635.204p 0 635.205p 10000.0u 635.206p 0 636.932p 0 636.933p 10000.0u 636.934p 0 642.902p 0 642.903p 10000.0u 642.904p 0 645.995p 0 645.996p 10000.0u 645.997p 0 651.479p 0 651.48p 10000.0u 651.481p 0 663.563p 0 663.564p 10000.0u 663.565p 0 674.291p 0 674.292p 10000.0u 674.293p 0 677.516p 0 677.517p 10000.0u 677.518p 0 679.115p 0 679.116p 10000.0u 679.117p 0 682.892p 0 682.893p 10000.0u 682.894p 0 685.106p 0 685.107p 10000.0u 685.108p 0 687.791p 0 687.792p 10000.0u 687.793p 0 710.924p 0 710.925p 10000.0u 710.926p 0 712.112p 0 712.113p 10000.0u 712.114p 0 747.107p 0 747.108p 10000.0u 747.109p 0 747.791p 0 747.792p 10000.0u 747.793p 0 748.52p 0 748.521p 10000.0u 748.522p 0 749.195p 0 749.196p 10000.0u 749.197p 0 750.23p 0 750.231p 10000.0u 750.232p 0 763.523p 0 763.524p 10000.0u 763.525p 0 769.286p 0 769.287p 10000.0u 769.288p 0 772.223p 0 772.224p 10000.0u 772.225p 0 813.125p 0 813.126p 10000.0u 813.127p 0 815.237p 0 815.238p 10000.0u 815.239p 0 817.19p 0 817.191p 10000.0u 817.192p 0 823.091p 0 823.092p 10000.0u 823.093p 0 827.42p 0 827.421p 10000.0u 827.422p 0 834.053p 0 834.054p 10000.0u 834.055p 0 846.767p 0 846.768p 10000.0u 846.769p 0 847.532p 0 847.533p 10000.0u 847.534p 0 869.726p 0 869.727p 10000.0u 869.728p 0 892.592p 0 892.593p 10000.0u 892.594p 0 911.414p 0 911.415p 10000.0u 911.416p 0 913.538p 0 913.539p 10000.0u 913.54p 0 923.897p 0 923.898p 10000.0u 923.899p 0 925.979p 0 925.98p 10000.0u 925.981p 0 943.991p 0 943.992p 10000.0u 943.993p 0 944.084p 0 944.085p 10000.0u 944.086p 0 945.38p 0 945.381p 10000.0u 945.382p 0 973.55p 0 973.551p 10000.0u 973.552p 0 977.813p 0 977.814p 10000.0u 977.815p 0 979.889p 0 979.89p 10000.0u 979.891p 0)
IIN36 0 37 pwl(0 0 2.984p 0 2.985p 10000.0u 2.986p 0 8.711p 0 8.712p 10000.0u 8.713p 0 19.91p 0 19.911p 10000.0u 19.912p 0 56.42p 0 56.421p 10000.0u 56.422p 0 58.229p 0 58.23p 10000.0u 58.231p 0 62.324p 0 62.325p 10000.0u 62.326p 0 65.153p 0 65.154p 10000.0u 65.155p 0 71.912p 0 71.913p 10000.0u 71.914p 0 74.942p 0 74.943p 10000.0u 74.944p 0 78.644p 0 78.645p 10000.0u 78.646p 0 81.812p 0 81.813p 10000.0u 81.814p 0 96.473p 0 96.474p 10000.0u 96.475p 0 102.62p 0 102.621p 10000.0u 102.622p 0 106.922p 0 106.923p 10000.0u 106.924p 0 117.656p 0 117.657p 10000.0u 117.658p 0 119.876p 0 119.877p 10000.0u 119.878p 0 123.683p 0 123.684p 10000.0u 123.685p 0 127.685p 0 127.686p 10000.0u 127.687p 0 128.795p 0 128.796p 10000.0u 128.797p 0 134.87p 0 134.871p 10000.0u 134.872p 0 157.787p 0 157.788p 10000.0u 157.789p 0 172.505p 0 172.506p 10000.0u 172.507p 0 177.32p 0 177.321p 10000.0u 177.322p 0 188.264p 0 188.265p 10000.0u 188.266p 0 191.309p 0 191.31p 10000.0u 191.311p 0 195.977p 0 195.978p 10000.0u 195.979p 0 209.54p 0 209.541p 10000.0u 209.542p 0 213.797p 0 213.798p 10000.0u 213.799p 0 234.89p 0 234.891p 10000.0u 234.892p 0 254.015p 0 254.016p 10000.0u 254.017p 0 255.248p 0 255.249p 10000.0u 255.25p 0 262.454p 0 262.455p 10000.0u 262.456p 0 263.729p 0 263.73p 10000.0u 263.731p 0 281.756p 0 281.757p 10000.0u 281.758p 0 320.747p 0 320.748p 10000.0u 320.749p 0 330.395p 0 330.396p 10000.0u 330.397p 0 340.838p 0 340.839p 10000.0u 340.84p 0 341.561p 0 341.562p 10000.0u 341.563p 0 346.175p 0 346.176p 10000.0u 346.177p 0 347.291p 0 347.292p 10000.0u 347.293p 0 352.649p 0 352.65p 10000.0u 352.651p 0 376.547p 0 376.548p 10000.0u 376.549p 0 377.456p 0 377.457p 10000.0u 377.458p 0 381.824p 0 381.825p 10000.0u 381.826p 0 384.896p 0 384.897p 10000.0u 384.898p 0 405.515p 0 405.516p 10000.0u 405.517p 0 412.346p 0 412.347p 10000.0u 412.348p 0 422.438p 0 422.439p 10000.0u 422.44p 0 436.772p 0 436.773p 10000.0u 436.774p 0 442.064p 0 442.065p 10000.0u 442.066p 0 442.721p 0 442.722p 10000.0u 442.723p 0 448.151p 0 448.152p 10000.0u 448.153p 0 465.926p 0 465.927p 10000.0u 465.928p 0 480.347p 0 480.348p 10000.0u 480.349p 0 481.316p 0 481.317p 10000.0u 481.318p 0 481.682p 0 481.683p 10000.0u 481.684p 0 482.327p 0 482.328p 10000.0u 482.329p 0 485.411p 0 485.412p 10000.0u 485.413p 0 488.027p 0 488.028p 10000.0u 488.029p 0 503.525p 0 503.526p 10000.0u 503.527p 0 510.431p 0 510.432p 10000.0u 510.433p 0 534.503p 0 534.504p 10000.0u 534.505p 0 545.003p 0 545.004p 10000.0u 545.005p 0 545.753p 0 545.754p 10000.0u 545.755p 0 560.09p 0 560.091p 10000.0u 560.092p 0 560.351p 0 560.352p 10000.0u 560.353p 0 566.549p 0 566.55p 10000.0u 566.551p 0 571.064p 0 571.065p 10000.0u 571.066p 0 574.991p 0 574.992p 10000.0u 574.993p 0 582.935p 0 582.936p 10000.0u 582.937p 0 586.16p 0 586.161p 10000.0u 586.162p 0 612.785p 0 612.786p 10000.0u 612.787p 0 627.188p 0 627.189p 10000.0u 627.19p 0 639.107p 0 639.108p 10000.0u 639.109p 0 643.298p 0 643.299p 10000.0u 643.3p 0 648.428p 0 648.429p 10000.0u 648.43p 0 650.465p 0 650.466p 10000.0u 650.467p 0 663.239p 0 663.24p 10000.0u 663.241p 0 682.679p 0 682.68p 10000.0u 682.681p 0 710.471p 0 710.472p 10000.0u 710.473p 0 724.514p 0 724.515p 10000.0u 724.516p 0 739.328p 0 739.329p 10000.0u 739.33p 0 749.708p 0 749.709p 10000.0u 749.71p 0 759.992p 0 759.993p 10000.0u 759.994p 0 763.433p 0 763.434p 10000.0u 763.435p 0 768.296p 0 768.297p 10000.0u 768.298p 0 777.956p 0 777.957p 10000.0u 777.958p 0 794.534p 0 794.535p 10000.0u 794.536p 0 799.13p 0 799.131p 10000.0u 799.132p 0 805.229p 0 805.23p 10000.0u 805.231p 0 834.422p 0 834.423p 10000.0u 834.424p 0 850.892p 0 850.893p 10000.0u 850.894p 0 861.83p 0 861.831p 10000.0u 861.832p 0 865.085p 0 865.086p 10000.0u 865.087p 0 898.481p 0 898.482p 10000.0u 898.483p 0 909.077p 0 909.078p 10000.0u 909.079p 0 911.843p 0 911.844p 10000.0u 911.845p 0 913.913p 0 913.914p 10000.0u 913.915p 0 914.45p 0 914.451p 10000.0u 914.452p 0 932.735p 0 932.736p 10000.0u 932.737p 0 945.176p 0 945.177p 10000.0u 945.178p 0 962.579p 0 962.58p 10000.0u 962.581p 0 974.369p 0 974.37p 10000.0u 974.371p 0 974.798p 0 974.799p 10000.0u 974.8p 0 982.676p 0 982.677p 10000.0u 982.678p 0)
IIN37 0 38 pwl(0 0 10.367p 0 10.368p 10000.0u 10.369p 0 28.256p 0 28.257p 10000.0u 28.258p 0 36.431p 0 36.432p 10000.0u 36.433p 0 59.879p 0 59.88p 10000.0u 59.881p 0 60.701p 0 60.702p 10000.0u 60.703p 0 83.483p 0 83.484p 10000.0u 83.485p 0 93.851p 0 93.852p 10000.0u 93.853p 0 102.314p 0 102.315p 10000.0u 102.316p 0 114.443p 0 114.444p 10000.0u 114.445p 0 125.561p 0 125.562p 10000.0u 125.563p 0 126.641p 0 126.642p 10000.0u 126.643p 0 146.933p 0 146.934p 10000.0u 146.935p 0 152.594p 0 152.595p 10000.0u 152.596p 0 159.14p 0 159.141p 10000.0u 159.142p 0 163.355p 0 163.356p 10000.0u 163.357p 0 165.902p 0 165.903p 10000.0u 165.904p 0 167.15p 0 167.151p 10000.0u 167.152p 0 167.744p 0 167.745p 10000.0u 167.746p 0 176.222p 0 176.223p 10000.0u 176.224p 0 177.26p 0 177.261p 10000.0u 177.262p 0 181.226p 0 181.227p 10000.0u 181.228p 0 184.535p 0 184.536p 10000.0u 184.537p 0 203.126p 0 203.127p 10000.0u 203.128p 0 208.007p 0 208.008p 10000.0u 208.009p 0 224.105p 0 224.106p 10000.0u 224.107p 0 240.014p 0 240.015p 10000.0u 240.016p 0 269.273p 0 269.274p 10000.0u 269.275p 0 270.107p 0 270.108p 10000.0u 270.109p 0 271.07p 0 271.071p 10000.0u 271.072p 0 284.813p 0 284.814p 10000.0u 284.815p 0 288.956p 0 288.957p 10000.0u 288.958p 0 293.549p 0 293.55p 10000.0u 293.551p 0 299.774p 0 299.775p 10000.0u 299.776p 0 310.517p 0 310.518p 10000.0u 310.519p 0 315.485p 0 315.486p 10000.0u 315.487p 0 322.271p 0 322.272p 10000.0u 322.273p 0 327.11p 0 327.111p 10000.0u 327.112p 0 328.508p 0 328.509p 10000.0u 328.51p 0 328.916p 0 328.917p 10000.0u 328.918p 0 354.062p 0 354.063p 10000.0u 354.064p 0 356.324p 0 356.325p 10000.0u 356.326p 0 357.269p 0 357.27p 10000.0u 357.271p 0 357.776p 0 357.777p 10000.0u 357.778p 0 368.654p 0 368.655p 10000.0u 368.656p 0 373.598p 0 373.599p 10000.0u 373.6p 0 398.588p 0 398.589p 10000.0u 398.59p 0 399.485p 0 399.486p 10000.0u 399.487p 0 413.351p 0 413.352p 10000.0u 413.353p 0 428.597p 0 428.598p 10000.0u 428.599p 0 441.869p 0 441.87p 10000.0u 441.871p 0 450.851p 0 450.852p 10000.0u 450.853p 0 459.641p 0 459.642p 10000.0u 459.643p 0 464.381p 0 464.382p 10000.0u 464.383p 0 465.206p 0 465.207p 10000.0u 465.208p 0 467.807p 0 467.808p 10000.0u 467.809p 0 491.141p 0 491.142p 10000.0u 491.143p 0 525.308p 0 525.309p 10000.0u 525.31p 0 525.527p 0 525.528p 10000.0u 525.529p 0 536.084p 0 536.085p 10000.0u 536.086p 0 554.228p 0 554.229p 10000.0u 554.23p 0 555.974p 0 555.975p 10000.0u 555.976p 0 571.751p 0 571.752p 10000.0u 571.753p 0 587.573p 0 587.574p 10000.0u 587.575p 0 593.501p 0 593.502p 10000.0u 593.503p 0 599.078p 0 599.079p 10000.0u 599.08p 0 605.153p 0 605.154p 10000.0u 605.155p 0 605.525p 0 605.526p 10000.0u 605.527p 0 616.547p 0 616.548p 10000.0u 616.549p 0 631.799p 0 631.8p 10000.0u 631.801p 0 633.536p 0 633.537p 10000.0u 633.538p 0 640.538p 0 640.539p 10000.0u 640.54p 0 684.038p 0 684.039p 10000.0u 684.04p 0 689.675p 0 689.676p 10000.0u 689.677p 0 698.231p 0 698.232p 10000.0u 698.233p 0 703.709p 0 703.71p 10000.0u 703.711p 0 715.43p 0 715.431p 10000.0u 715.432p 0 735.164p 0 735.165p 10000.0u 735.166p 0 764.528p 0 764.529p 10000.0u 764.53p 0 777.026p 0 777.027p 10000.0u 777.028p 0 778.157p 0 778.158p 10000.0u 778.159p 0 784.754p 0 784.755p 10000.0u 784.756p 0 802.379p 0 802.38p 10000.0u 802.381p 0 844.154p 0 844.155p 10000.0u 844.156p 0 865.223p 0 865.224p 10000.0u 865.225p 0 866.912p 0 866.913p 10000.0u 866.914p 0 890.444p 0 890.445p 10000.0u 890.446p 0 896.345p 0 896.346p 10000.0u 896.347p 0 900.2p 0 900.201p 10000.0u 900.202p 0 930.542p 0 930.543p 10000.0u 930.544p 0 937.454p 0 937.455p 10000.0u 937.456p 0 938.879p 0 938.88p 10000.0u 938.881p 0 942.254p 0 942.255p 10000.0u 942.256p 0 946.694p 0 946.695p 10000.0u 946.696p 0 952.577p 0 952.578p 10000.0u 952.579p 0 962.132p 0 962.133p 10000.0u 962.134p 0 970.955p 0 970.956p 10000.0u 970.957p 0 974.387p 0 974.388p 10000.0u 974.389p 0 976.01p 0 976.011p 10000.0u 976.012p 0 997.088p 0 997.089p 10000.0u 997.09p 0)
IIN38 0 39 pwl(0 0 2.369p 0 2.37p 10000.0u 2.371p 0 15.617p 0 15.618p 10000.0u 15.619p 0 15.98p 0 15.981p 10000.0u 15.982p 0 38.009p 0 38.01p 10000.0u 38.011p 0 50.3p 0 50.301p 10000.0u 50.302p 0 59.399p 0 59.4p 10000.0u 59.401p 0 68.786p 0 68.787p 10000.0u 68.788p 0 78.008p 0 78.009p 10000.0u 78.01p 0 83.837p 0 83.838p 10000.0u 83.839p 0 129.818p 0 129.819p 10000.0u 129.82p 0 135.743p 0 135.744p 10000.0u 135.745p 0 149.936p 0 149.937p 10000.0u 149.938p 0 155.453p 0 155.454p 10000.0u 155.455p 0 164.63p 0 164.631p 10000.0u 164.632p 0 175.013p 0 175.014p 10000.0u 175.015p 0 186.251p 0 186.252p 10000.0u 186.253p 0 187.229p 0 187.23p 10000.0u 187.231p 0 212.933p 0 212.934p 10000.0u 212.935p 0 218.354p 0 218.355p 10000.0u 218.356p 0 235.412p 0 235.413p 10000.0u 235.414p 0 295.991p 0 295.992p 10000.0u 295.993p 0 315.71p 0 315.711p 10000.0u 315.712p 0 322.316p 0 322.317p 10000.0u 322.318p 0 326.213p 0 326.214p 10000.0u 326.215p 0 332.957p 0 332.958p 10000.0u 332.959p 0 335.447p 0 335.448p 10000.0u 335.449p 0 338.576p 0 338.577p 10000.0u 338.578p 0 363.047p 0 363.048p 10000.0u 363.049p 0 365.525p 0 365.526p 10000.0u 365.527p 0 366.32p 0 366.321p 10000.0u 366.322p 0 367.733p 0 367.734p 10000.0u 367.735p 0 372.932p 0 372.933p 10000.0u 372.934p 0 375.29p 0 375.291p 10000.0u 375.292p 0 380.555p 0 380.556p 10000.0u 380.557p 0 399.365p 0 399.366p 10000.0u 399.367p 0 413.753p 0 413.754p 10000.0u 413.755p 0 442.337p 0 442.338p 10000.0u 442.339p 0 443.504p 0 443.505p 10000.0u 443.506p 0 445.388p 0 445.389p 10000.0u 445.39p 0 463.31p 0 463.311p 10000.0u 463.312p 0 482.303p 0 482.304p 10000.0u 482.305p 0 518.786p 0 518.787p 10000.0u 518.788p 0 529.211p 0 529.212p 10000.0u 529.213p 0 541.793p 0 541.794p 10000.0u 541.795p 0 543.116p 0 543.117p 10000.0u 543.118p 0 550.196p 0 550.197p 10000.0u 550.198p 0 559.397p 0 559.398p 10000.0u 559.399p 0 560.51p 0 560.511p 10000.0u 560.512p 0 570.725p 0 570.726p 10000.0u 570.727p 0 571.988p 0 571.989p 10000.0u 571.99p 0 596.327p 0 596.328p 10000.0u 596.329p 0 597.668p 0 597.669p 10000.0u 597.67p 0 641.828p 0 641.829p 10000.0u 641.83p 0 645.683p 0 645.684p 10000.0u 645.685p 0 648.278p 0 648.279p 10000.0u 648.28p 0 650.198p 0 650.199p 10000.0u 650.2p 0 655.625p 0 655.626p 10000.0u 655.627p 0 655.949p 0 655.95p 10000.0u 655.951p 0 656.39p 0 656.391p 10000.0u 656.392p 0 676.19p 0 676.191p 10000.0u 676.192p 0 685.511p 0 685.512p 10000.0u 685.513p 0 716.759p 0 716.76p 10000.0u 716.761p 0 737.228p 0 737.229p 10000.0u 737.23p 0 767.882p 0 767.883p 10000.0u 767.884p 0 790.142p 0 790.143p 10000.0u 790.144p 0 800.714p 0 800.715p 10000.0u 800.716p 0 815.828p 0 815.829p 10000.0u 815.83p 0 818.447p 0 818.448p 10000.0u 818.449p 0 820.673p 0 820.674p 10000.0u 820.675p 0 845.477p 0 845.478p 10000.0u 845.479p 0 851.882p 0 851.883p 10000.0u 851.884p 0 862.22p 0 862.221p 10000.0u 862.222p 0 890.15p 0 890.151p 10000.0u 890.152p 0 892.247p 0 892.248p 10000.0u 892.249p 0 929.342p 0 929.343p 10000.0u 929.344p 0 966.383p 0 966.384p 10000.0u 966.385p 0 971.582p 0 971.583p 10000.0u 971.584p 0)
IIN39 0 40 pwl(0 0 4.019p 0 4.02p 10000.0u 4.021p 0 36.896p 0 36.897p 10000.0u 36.898p 0 38.759p 0 38.76p 10000.0u 38.761p 0 46.934p 0 46.935p 10000.0u 46.936p 0 59.903p 0 59.904p 10000.0u 59.905p 0 62.369p 0 62.37p 10000.0u 62.371p 0 76.193p 0 76.194p 10000.0u 76.195p 0 83.552p 0 83.553p 10000.0u 83.554p 0 91.028p 0 91.029p 10000.0u 91.03p 0 101.657p 0 101.658p 10000.0u 101.659p 0 111.44p 0 111.441p 10000.0u 111.442p 0 133.256p 0 133.257p 10000.0u 133.258p 0 147.701p 0 147.702p 10000.0u 147.703p 0 155.012p 0 155.013p 10000.0u 155.014p 0 156.305p 0 156.306p 10000.0u 156.307p 0 160.25p 0 160.251p 10000.0u 160.252p 0 165.311p 0 165.312p 10000.0u 165.313p 0 185.663p 0 185.664p 10000.0u 185.665p 0 190.451p 0 190.452p 10000.0u 190.453p 0 199.394p 0 199.395p 10000.0u 199.396p 0 206.666p 0 206.667p 10000.0u 206.668p 0 218.69p 0 218.691p 10000.0u 218.692p 0 227.72p 0 227.721p 10000.0u 227.722p 0 233.816p 0 233.817p 10000.0u 233.818p 0 258.023p 0 258.024p 10000.0u 258.025p 0 260.78p 0 260.781p 10000.0u 260.782p 0 264.554p 0 264.555p 10000.0u 264.556p 0 269.018p 0 269.019p 10000.0u 269.02p 0 270.491p 0 270.492p 10000.0u 270.493p 0 273.782p 0 273.783p 10000.0u 273.784p 0 299.978p 0 299.979p 10000.0u 299.98p 0 301.283p 0 301.284p 10000.0u 301.285p 0 337.232p 0 337.233p 10000.0u 337.234p 0 341.528p 0 341.529p 10000.0u 341.53p 0 349.301p 0 349.302p 10000.0u 349.303p 0 369.893p 0 369.894p 10000.0u 369.895p 0 371.042p 0 371.043p 10000.0u 371.044p 0 371.273p 0 371.274p 10000.0u 371.275p 0 393.809p 0 393.81p 10000.0u 393.811p 0 400.337p 0 400.338p 10000.0u 400.339p 0 403.364p 0 403.365p 10000.0u 403.366p 0 412.238p 0 412.239p 10000.0u 412.24p 0 433.118p 0 433.119p 10000.0u 433.12p 0 436.973p 0 436.974p 10000.0u 436.975p 0 437.849p 0 437.85p 10000.0u 437.851p 0 443.696p 0 443.697p 10000.0u 443.698p 0 445.382p 0 445.383p 10000.0u 445.384p 0 453.869p 0 453.87p 10000.0u 453.871p 0 488.036p 0 488.037p 10000.0u 488.038p 0 488.216p 0 488.217p 10000.0u 488.218p 0 497.723p 0 497.724p 10000.0u 497.725p 0 501.062p 0 501.063p 10000.0u 501.064p 0 524.282p 0 524.283p 10000.0u 524.284p 0 530.84p 0 530.841p 10000.0u 530.842p 0 548.408p 0 548.409p 10000.0u 548.41p 0 554.612p 0 554.613p 10000.0u 554.614p 0 555.539p 0 555.54p 10000.0u 555.541p 0 569.858p 0 569.859p 10000.0u 569.86p 0 572.624p 0 572.625p 10000.0u 572.626p 0 575.627p 0 575.628p 10000.0u 575.629p 0 578.204p 0 578.205p 10000.0u 578.206p 0 588.131p 0 588.132p 10000.0u 588.133p 0 598.502p 0 598.503p 10000.0u 598.504p 0 613.28p 0 613.281p 10000.0u 613.282p 0 621.764p 0 621.765p 10000.0u 621.766p 0 629.024p 0 629.025p 10000.0u 629.026p 0 630.968p 0 630.969p 10000.0u 630.97p 0 647.312p 0 647.313p 10000.0u 647.314p 0 664.973p 0 664.974p 10000.0u 664.975p 0 667.613p 0 667.614p 10000.0u 667.615p 0 678.62p 0 678.621p 10000.0u 678.622p 0 682.553p 0 682.554p 10000.0u 682.555p 0 682.928p 0 682.929p 10000.0u 682.93p 0 700.829p 0 700.83p 10000.0u 700.831p 0 706.1p 0 706.101p 10000.0u 706.102p 0 720.38p 0 720.381p 10000.0u 720.382p 0 738.761p 0 738.762p 10000.0u 738.763p 0 742.349p 0 742.35p 10000.0u 742.351p 0 767.018p 0 767.019p 10000.0u 767.02p 0 772.028p 0 772.029p 10000.0u 772.03p 0 772.442p 0 772.443p 10000.0u 772.444p 0 775.595p 0 775.596p 10000.0u 775.597p 0 778.022p 0 778.023p 10000.0u 778.024p 0 784.61p 0 784.611p 10000.0u 784.612p 0 784.691p 0 784.692p 10000.0u 784.693p 0 786.152p 0 786.153p 10000.0u 786.154p 0 789.347p 0 789.348p 10000.0u 789.349p 0 794.258p 0 794.259p 10000.0u 794.26p 0 796.247p 0 796.248p 10000.0u 796.249p 0 802.712p 0 802.713p 10000.0u 802.714p 0 803.927p 0 803.928p 10000.0u 803.929p 0 806.906p 0 806.907p 10000.0u 806.908p 0 810.05p 0 810.051p 10000.0u 810.052p 0 811.358p 0 811.359p 10000.0u 811.36p 0 811.898p 0 811.899p 10000.0u 811.9p 0 815.774p 0 815.775p 10000.0u 815.776p 0 815.783p 0 815.784p 10000.0u 815.785p 0 817.073p 0 817.074p 10000.0u 817.075p 0 818.156p 0 818.157p 10000.0u 818.158p 0 833.585p 0 833.586p 10000.0u 833.587p 0 836.786p 0 836.787p 10000.0u 836.788p 0 839.9p 0 839.901p 10000.0u 839.902p 0 857.066p 0 857.067p 10000.0u 857.068p 0 857.831p 0 857.832p 10000.0u 857.833p 0 862.103p 0 862.104p 10000.0u 862.105p 0 877.55p 0 877.551p 10000.0u 877.552p 0 885.95p 0 885.951p 10000.0u 885.952p 0 892.505p 0 892.506p 10000.0u 892.507p 0 893.294p 0 893.295p 10000.0u 893.296p 0 923.516p 0 923.517p 10000.0u 923.518p 0 944.54p 0 944.541p 10000.0u 944.542p 0 951.047p 0 951.048p 10000.0u 951.049p 0 951.707p 0 951.708p 10000.0u 951.709p 0 952.436p 0 952.437p 10000.0u 952.438p 0 956.612p 0 956.613p 10000.0u 956.614p 0 966.236p 0 966.237p 10000.0u 966.238p 0 970.169p 0 970.17p 10000.0u 970.171p 0)
IIN40 0 41 pwl(0 0 2.585p 0 2.586p 10000.0u 2.587p 0 19.316p 0 19.317p 10000.0u 19.318p 0 42.812p 0 42.813p 10000.0u 42.814p 0 48.599p 0 48.6p 10000.0u 48.601p 0 55.469p 0 55.47p 10000.0u 55.471p 0 63.854p 0 63.855p 10000.0u 63.856p 0 72.26p 0 72.261p 10000.0u 72.262p 0 93.857p 0 93.858p 10000.0u 93.859p 0 100.148p 0 100.149p 10000.0u 100.15p 0 124.205p 0 124.206p 10000.0u 124.207p 0 130.115p 0 130.116p 10000.0u 130.117p 0 130.514p 0 130.515p 10000.0u 130.516p 0 143.963p 0 143.964p 10000.0u 143.965p 0 150.671p 0 150.672p 10000.0u 150.673p 0 172.103p 0 172.104p 10000.0u 172.105p 0 180.317p 0 180.318p 10000.0u 180.319p 0 192.542p 0 192.543p 10000.0u 192.544p 0 198.536p 0 198.537p 10000.0u 198.538p 0 208.277p 0 208.278p 10000.0u 208.279p 0 218.342p 0 218.343p 10000.0u 218.344p 0 220.145p 0 220.146p 10000.0u 220.147p 0 232.436p 0 232.437p 10000.0u 232.438p 0 232.946p 0 232.947p 10000.0u 232.948p 0 233.477p 0 233.478p 10000.0u 233.479p 0 234.614p 0 234.615p 10000.0u 234.616p 0 238.991p 0 238.992p 10000.0u 238.993p 0 240.602p 0 240.603p 10000.0u 240.604p 0 242.699p 0 242.7p 10000.0u 242.701p 0 242.819p 0 242.82p 10000.0u 242.821p 0 254.021p 0 254.022p 10000.0u 254.023p 0 259.715p 0 259.716p 10000.0u 259.717p 0 261.641p 0 261.642p 10000.0u 261.643p 0 263.738p 0 263.739p 10000.0u 263.74p 0 284.987p 0 284.988p 10000.0u 284.989p 0 305.579p 0 305.58p 10000.0u 305.581p 0 311.846p 0 311.847p 10000.0u 311.848p 0 317.327p 0 317.328p 10000.0u 317.329p 0 344.321p 0 344.322p 10000.0u 344.323p 0 352.955p 0 352.956p 10000.0u 352.957p 0 356.966p 0 356.967p 10000.0u 356.968p 0 364.802p 0 364.803p 10000.0u 364.804p 0 381.836p 0 381.837p 10000.0u 381.838p 0 382.79p 0 382.791p 10000.0u 382.792p 0 389.549p 0 389.55p 10000.0u 389.551p 0 391.982p 0 391.983p 10000.0u 391.984p 0 398.294p 0 398.295p 10000.0u 398.296p 0 406.481p 0 406.482p 10000.0u 406.483p 0 427.271p 0 427.272p 10000.0u 427.273p 0 427.535p 0 427.536p 10000.0u 427.537p 0 439.991p 0 439.992p 10000.0u 439.993p 0 482.546p 0 482.547p 10000.0u 482.548p 0 484.487p 0 484.488p 10000.0u 484.489p 0 487.505p 0 487.506p 10000.0u 487.507p 0 496.274p 0 496.275p 10000.0u 496.276p 0 503.588p 0 503.589p 10000.0u 503.59p 0 505.211p 0 505.212p 10000.0u 505.213p 0 522.137p 0 522.138p 10000.0u 522.139p 0 528.968p 0 528.969p 10000.0u 528.97p 0 539.381p 0 539.382p 10000.0u 539.383p 0 557.243p 0 557.244p 10000.0u 557.245p 0 563.792p 0 563.793p 10000.0u 563.794p 0 585.05p 0 585.051p 10000.0u 585.052p 0 586.988p 0 586.989p 10000.0u 586.99p 0 589.217p 0 589.218p 10000.0u 589.219p 0 605.474p 0 605.475p 10000.0u 605.476p 0 612.305p 0 612.306p 10000.0u 612.307p 0 620.864p 0 620.865p 10000.0u 620.866p 0 622.103p 0 622.104p 10000.0u 622.105p 0 623.351p 0 623.352p 10000.0u 623.353p 0 630.077p 0 630.078p 10000.0u 630.079p 0 632.522p 0 632.523p 10000.0u 632.524p 0 638.975p 0 638.976p 10000.0u 638.977p 0 662.369p 0 662.37p 10000.0u 662.371p 0 684.812p 0 684.813p 10000.0u 684.814p 0 712.217p 0 712.218p 10000.0u 712.219p 0 713.516p 0 713.517p 10000.0u 713.518p 0 715.418p 0 715.419p 10000.0u 715.42p 0 724.979p 0 724.98p 10000.0u 724.981p 0 727.925p 0 727.926p 10000.0u 727.927p 0 743.54p 0 743.541p 10000.0u 743.542p 0 766.529p 0 766.53p 10000.0u 766.531p 0 817.229p 0 817.23p 10000.0u 817.231p 0 823.535p 0 823.536p 10000.0u 823.537p 0 832.391p 0 832.392p 10000.0u 832.393p 0 833.102p 0 833.103p 10000.0u 833.104p 0 833.387p 0 833.388p 10000.0u 833.389p 0 868.862p 0 868.863p 10000.0u 868.864p 0 874.583p 0 874.584p 10000.0u 874.585p 0 889.478p 0 889.479p 10000.0u 889.48p 0 897.434p 0 897.435p 10000.0u 897.436p 0 907.181p 0 907.182p 10000.0u 907.183p 0 924.134p 0 924.135p 10000.0u 924.136p 0 924.458p 0 924.459p 10000.0u 924.46p 0 927.479p 0 927.48p 10000.0u 927.481p 0 931.838p 0 931.839p 10000.0u 931.84p 0 939.398p 0 939.399p 10000.0u 939.4p 0 942.716p 0 942.717p 10000.0u 942.718p 0 942.92p 0 942.921p 10000.0u 942.922p 0 952.178p 0 952.179p 10000.0u 952.18p 0 964.532p 0 964.533p 10000.0u 964.534p 0 965.126p 0 965.127p 10000.0u 965.128p 0 965.861p 0 965.862p 10000.0u 965.863p 0 973.559p 0 973.56p 10000.0u 973.561p 0 988.961p 0 988.962p 10000.0u 988.963p 0 991.475p 0 991.476p 10000.0u 991.477p 0)
IIN41 0 42 pwl(0 0 2.747p 0 2.748p 10000.0u 2.749p 0 3.893p 0 3.894p 10000.0u 3.895p 0 6.125p 0 6.126p 10000.0u 6.127p 0 18.956p 0 18.957p 10000.0u 18.958p 0 23.612p 0 23.613p 10000.0u 23.614p 0 34.427p 0 34.428p 10000.0u 34.429p 0 43.22p 0 43.221p 10000.0u 43.222p 0 62.354p 0 62.355p 10000.0u 62.356p 0 68.903p 0 68.904p 10000.0u 68.905p 0 82.574p 0 82.575p 10000.0u 82.576p 0 92.855p 0 92.856p 10000.0u 92.857p 0 93.596p 0 93.597p 10000.0u 93.598p 0 106.634p 0 106.635p 10000.0u 106.636p 0 117.686p 0 117.687p 10000.0u 117.688p 0 121.361p 0 121.362p 10000.0u 121.363p 0 131.819p 0 131.82p 10000.0u 131.821p 0 132.068p 0 132.069p 10000.0u 132.07p 0 152.972p 0 152.973p 10000.0u 152.974p 0 175.223p 0 175.224p 10000.0u 175.225p 0 191.594p 0 191.595p 10000.0u 191.596p 0 194.426p 0 194.427p 10000.0u 194.428p 0 194.63p 0 194.631p 10000.0u 194.632p 0 202.52p 0 202.521p 10000.0u 202.522p 0 204.179p 0 204.18p 10000.0u 204.181p 0 220.712p 0 220.713p 10000.0u 220.714p 0 227.33p 0 227.331p 10000.0u 227.332p 0 232.355p 0 232.356p 10000.0u 232.357p 0 276.965p 0 276.966p 10000.0u 276.967p 0 277.946p 0 277.947p 10000.0u 277.948p 0 284.996p 0 284.997p 10000.0u 284.998p 0 285.884p 0 285.885p 10000.0u 285.886p 0 299.687p 0 299.688p 10000.0u 299.689p 0 302.9p 0 302.901p 10000.0u 302.902p 0 303.599p 0 303.6p 10000.0u 303.601p 0 320.546p 0 320.547p 10000.0u 320.548p 0 333.704p 0 333.705p 10000.0u 333.706p 0 362.3p 0 362.301p 10000.0u 362.302p 0 364.592p 0 364.593p 10000.0u 364.594p 0 385.106p 0 385.107p 10000.0u 385.108p 0 390.257p 0 390.258p 10000.0u 390.259p 0 390.59p 0 390.591p 10000.0u 390.592p 0 397.682p 0 397.683p 10000.0u 397.684p 0 438.107p 0 438.108p 10000.0u 438.109p 0 444.305p 0 444.306p 10000.0u 444.307p 0 444.899p 0 444.9p 10000.0u 444.901p 0 455.858p 0 455.859p 10000.0u 455.86p 0 456.806p 0 456.807p 10000.0u 456.808p 0 466.304p 0 466.305p 10000.0u 466.306p 0 473.078p 0 473.079p 10000.0u 473.08p 0 474.578p 0 474.579p 10000.0u 474.58p 0 477.752p 0 477.753p 10000.0u 477.754p 0 479.306p 0 479.307p 10000.0u 479.308p 0 490.937p 0 490.938p 10000.0u 490.939p 0 493.76p 0 493.761p 10000.0u 493.762p 0 502.553p 0 502.554p 10000.0u 502.555p 0 504.242p 0 504.243p 10000.0u 504.244p 0 511.226p 0 511.227p 10000.0u 511.228p 0 514.118p 0 514.119p 10000.0u 514.12p 0 515.21p 0 515.211p 10000.0u 515.212p 0 530.855p 0 530.856p 10000.0u 530.857p 0 548.432p 0 548.433p 10000.0u 548.434p 0 549.782p 0 549.783p 10000.0u 549.784p 0 563.003p 0 563.004p 10000.0u 563.005p 0 564.593p 0 564.594p 10000.0u 564.595p 0 566.105p 0 566.106p 10000.0u 566.107p 0 566.546p 0 566.547p 10000.0u 566.548p 0 574.298p 0 574.299p 10000.0u 574.3p 0 593.801p 0 593.802p 10000.0u 593.803p 0 620.525p 0 620.526p 10000.0u 620.527p 0 632.948p 0 632.949p 10000.0u 632.95p 0 636.875p 0 636.876p 10000.0u 636.877p 0 648.344p 0 648.345p 10000.0u 648.346p 0 656.288p 0 656.289p 10000.0u 656.29p 0 673.775p 0 673.776p 10000.0u 673.777p 0 728.84p 0 728.841p 10000.0u 728.842p 0 778.298p 0 778.299p 10000.0u 778.3p 0 779.726p 0 779.727p 10000.0u 779.728p 0 779.906p 0 779.907p 10000.0u 779.908p 0 783.323p 0 783.324p 10000.0u 783.325p 0 783.59p 0 783.591p 10000.0u 783.592p 0 851.699p 0 851.7p 10000.0u 851.701p 0 854.078p 0 854.079p 10000.0u 854.08p 0 882.545p 0 882.546p 10000.0u 882.547p 0 883.673p 0 883.674p 10000.0u 883.675p 0 917.756p 0 917.757p 10000.0u 917.758p 0 930.437p 0 930.438p 10000.0u 930.439p 0 932.12p 0 932.121p 10000.0u 932.122p 0 935.261p 0 935.262p 10000.0u 935.263p 0 967.823p 0 967.824p 10000.0u 967.825p 0 977.468p 0 977.469p 10000.0u 977.47p 0 993.626p 0 993.627p 10000.0u 993.628p 0 998.435p 0 998.436p 10000.0u 998.437p 0)
IIN42 0 43 pwl(0 0 11.792p 0 11.793p 10000.0u 11.794p 0 14.498p 0 14.499p 10000.0u 14.5p 0 21.32p 0 21.321p 10000.0u 21.322p 0 24.065p 0 24.066p 10000.0u 24.067p 0 28.244p 0 28.245p 10000.0u 28.246p 0 28.565p 0 28.566p 10000.0u 28.567p 0 31.769p 0 31.77p 10000.0u 31.771p 0 40.151p 0 40.152p 10000.0u 40.153p 0 50.582p 0 50.583p 10000.0u 50.584p 0 66.326p 0 66.327p 10000.0u 66.328p 0 69.596p 0 69.597p 10000.0u 69.598p 0 84.17p 0 84.171p 10000.0u 84.172p 0 85.262p 0 85.263p 10000.0u 85.264p 0 101.285p 0 101.286p 10000.0u 101.287p 0 110.267p 0 110.268p 10000.0u 110.269p 0 122.642p 0 122.643p 10000.0u 122.644p 0 126.443p 0 126.444p 10000.0u 126.445p 0 127.562p 0 127.563p 10000.0u 127.564p 0 133.916p 0 133.917p 10000.0u 133.918p 0 173.615p 0 173.616p 10000.0u 173.617p 0 177.575p 0 177.576p 10000.0u 177.577p 0 190.919p 0 190.92p 10000.0u 190.921p 0 200.186p 0 200.187p 10000.0u 200.188p 0 213.29p 0 213.291p 10000.0u 213.292p 0 230.711p 0 230.712p 10000.0u 230.713p 0 239.3p 0 239.301p 10000.0u 239.302p 0 247.853p 0 247.854p 10000.0u 247.855p 0 253.892p 0 253.893p 10000.0u 253.894p 0 265.349p 0 265.35p 10000.0u 265.351p 0 278.195p 0 278.196p 10000.0u 278.197p 0 283.964p 0 283.965p 10000.0u 283.966p 0 289.112p 0 289.113p 10000.0u 289.114p 0 300.41p 0 300.411p 10000.0u 300.412p 0 307.619p 0 307.62p 10000.0u 307.621p 0 325.772p 0 325.773p 10000.0u 325.774p 0 327.626p 0 327.627p 10000.0u 327.628p 0 329.288p 0 329.289p 10000.0u 329.29p 0 333.986p 0 333.987p 10000.0u 333.988p 0 334.805p 0 334.806p 10000.0u 334.807p 0 345.965p 0 345.966p 10000.0u 345.967p 0 347.243p 0 347.244p 10000.0u 347.245p 0 352.292p 0 352.293p 10000.0u 352.294p 0 363.14p 0 363.141p 10000.0u 363.142p 0 368.753p 0 368.754p 10000.0u 368.755p 0 396.44p 0 396.441p 10000.0u 396.442p 0 424.202p 0 424.203p 10000.0u 424.204p 0 425.651p 0 425.652p 10000.0u 425.653p 0 429.053p 0 429.054p 10000.0u 429.055p 0 437.078p 0 437.079p 10000.0u 437.08p 0 440.567p 0 440.568p 10000.0u 440.569p 0 453.179p 0 453.18p 10000.0u 453.181p 0 471.665p 0 471.666p 10000.0u 471.667p 0 474.512p 0 474.513p 10000.0u 474.514p 0 476.978p 0 476.979p 10000.0u 476.98p 0 505.694p 0 505.695p 10000.0u 505.696p 0 520.928p 0 520.929p 10000.0u 520.93p 0 554.531p 0 554.532p 10000.0u 554.533p 0 556.196p 0 556.197p 10000.0u 556.198p 0 567.074p 0 567.075p 10000.0u 567.076p 0 576.368p 0 576.369p 10000.0u 576.37p 0 596.057p 0 596.058p 10000.0u 596.059p 0 608.57p 0 608.571p 10000.0u 608.572p 0 609.431p 0 609.432p 10000.0u 609.433p 0 612.338p 0 612.339p 10000.0u 612.34p 0 623.183p 0 623.184p 10000.0u 623.185p 0 627.266p 0 627.267p 10000.0u 627.268p 0 629.291p 0 629.292p 10000.0u 629.293p 0 651.038p 0 651.039p 10000.0u 651.04p 0 663.956p 0 663.957p 10000.0u 663.958p 0 666.35p 0 666.351p 10000.0u 666.352p 0 671.549p 0 671.55p 10000.0u 671.551p 0 683.894p 0 683.895p 10000.0u 683.896p 0 686.447p 0 686.448p 10000.0u 686.449p 0 689.423p 0 689.424p 10000.0u 689.425p 0 691.286p 0 691.287p 10000.0u 691.288p 0 701.036p 0 701.037p 10000.0u 701.038p 0 713.786p 0 713.787p 10000.0u 713.788p 0 720.497p 0 720.498p 10000.0u 720.499p 0 729.998p 0 729.999p 10000.0u 730.0p 0 737.174p 0 737.175p 10000.0u 737.176p 0 738.953p 0 738.954p 10000.0u 738.955p 0 755.204p 0 755.205p 10000.0u 755.206p 0 758.57p 0 758.571p 10000.0u 758.572p 0 804.857p 0 804.858p 10000.0u 804.859p 0 814.367p 0 814.368p 10000.0u 814.369p 0 815.828p 0 815.829p 10000.0u 815.83p 0 824.429p 0 824.43p 10000.0u 824.431p 0 837.23p 0 837.231p 10000.0u 837.232p 0 840.389p 0 840.39p 10000.0u 840.391p 0 863.618p 0 863.619p 10000.0u 863.62p 0 871.889p 0 871.89p 10000.0u 871.891p 0 872.357p 0 872.358p 10000.0u 872.359p 0 890.96p 0 890.961p 10000.0u 890.962p 0 918.323p 0 918.324p 10000.0u 918.325p 0 929.873p 0 929.874p 10000.0u 929.875p 0 937.412p 0 937.413p 10000.0u 937.414p 0 945.983p 0 945.984p 10000.0u 945.985p 0 953.801p 0 953.802p 10000.0u 953.803p 0 963.38p 0 963.381p 10000.0u 963.382p 0 967.619p 0 967.62p 10000.0u 967.621p 0 985.226p 0 985.227p 10000.0u 985.228p 0)
IIN43 0 44 pwl(0 0 12.974p 0 12.975p 10000.0u 12.976p 0 15.185p 0 15.186p 10000.0u 15.187p 0 39.305p 0 39.306p 10000.0u 39.307p 0 41.087p 0 41.088p 10000.0u 41.089p 0 63.941p 0 63.942p 10000.0u 63.943p 0 67.52p 0 67.521p 10000.0u 67.522p 0 89.162p 0 89.163p 10000.0u 89.164p 0 94.88p 0 94.881p 10000.0u 94.882p 0 106.922p 0 106.923p 10000.0u 106.924p 0 117.743p 0 117.744p 10000.0u 117.745p 0 120.026p 0 120.027p 10000.0u 120.028p 0 124.925p 0 124.926p 10000.0u 124.927p 0 128.027p 0 128.028p 10000.0u 128.029p 0 162.449p 0 162.45p 10000.0u 162.451p 0 171.929p 0 171.93p 10000.0u 171.931p 0 177.398p 0 177.399p 10000.0u 177.4p 0 183.653p 0 183.654p 10000.0u 183.655p 0 186.767p 0 186.768p 10000.0u 186.769p 0 195.656p 0 195.657p 10000.0u 195.658p 0 205.571p 0 205.572p 10000.0u 205.573p 0 208.544p 0 208.545p 10000.0u 208.546p 0 215.645p 0 215.646p 10000.0u 215.647p 0 250.817p 0 250.818p 10000.0u 250.819p 0 250.892p 0 250.893p 10000.0u 250.894p 0 252.821p 0 252.822p 10000.0u 252.823p 0 264.074p 0 264.075p 10000.0u 264.076p 0 265.811p 0 265.812p 10000.0u 265.813p 0 266.504p 0 266.505p 10000.0u 266.506p 0 285.863p 0 285.864p 10000.0u 285.865p 0 307.502p 0 307.503p 10000.0u 307.504p 0 330.95p 0 330.951p 10000.0u 330.952p 0 331.412p 0 331.413p 10000.0u 331.414p 0 333.914p 0 333.915p 10000.0u 333.916p 0 340.838p 0 340.839p 10000.0u 340.84p 0 356.216p 0 356.217p 10000.0u 356.218p 0 367.454p 0 367.455p 10000.0u 367.456p 0 369.329p 0 369.33p 10000.0u 369.331p 0 397.814p 0 397.815p 10000.0u 397.816p 0 401.81p 0 401.811p 10000.0u 401.812p 0 429.113p 0 429.114p 10000.0u 429.115p 0 433.319p 0 433.32p 10000.0u 433.321p 0 435.998p 0 435.999p 10000.0u 436.0p 0 445.34p 0 445.341p 10000.0u 445.342p 0 451.292p 0 451.293p 10000.0u 451.294p 0 465.593p 0 465.594p 10000.0u 465.595p 0 484.322p 0 484.323p 10000.0u 484.324p 0 484.667p 0 484.668p 10000.0u 484.669p 0 492.896p 0 492.897p 10000.0u 492.898p 0 496.928p 0 496.929p 10000.0u 496.93p 0 498.479p 0 498.48p 10000.0u 498.481p 0 499.913p 0 499.914p 10000.0u 499.915p 0 528.428p 0 528.429p 10000.0u 528.43p 0 531.014p 0 531.015p 10000.0u 531.016p 0 556.178p 0 556.179p 10000.0u 556.18p 0 564.878p 0 564.879p 10000.0u 564.88p 0 568.208p 0 568.209p 10000.0u 568.21p 0 568.916p 0 568.917p 10000.0u 568.918p 0 569.849p 0 569.85p 10000.0u 569.851p 0 572.342p 0 572.343p 10000.0u 572.344p 0 577.154p 0 577.155p 10000.0u 577.156p 0 591.677p 0 591.678p 10000.0u 591.679p 0 606.809p 0 606.81p 10000.0u 606.811p 0 619.382p 0 619.383p 10000.0u 619.384p 0 622.979p 0 622.98p 10000.0u 622.981p 0 636.935p 0 636.936p 10000.0u 636.937p 0 639.083p 0 639.084p 10000.0u 639.085p 0 644.957p 0 644.958p 10000.0u 644.959p 0 646.184p 0 646.185p 10000.0u 646.186p 0 648.041p 0 648.042p 10000.0u 648.043p 0 660.59p 0 660.591p 10000.0u 660.592p 0 672.971p 0 672.972p 10000.0u 672.973p 0 692.822p 0 692.823p 10000.0u 692.824p 0 725.759p 0 725.76p 10000.0u 725.761p 0 736.925p 0 736.926p 10000.0u 736.927p 0 768.461p 0 768.462p 10000.0u 768.463p 0 769.838p 0 769.839p 10000.0u 769.84p 0 771.797p 0 771.798p 10000.0u 771.799p 0 775.127p 0 775.128p 10000.0u 775.129p 0 785.912p 0 785.913p 10000.0u 785.914p 0 792.164p 0 792.165p 10000.0u 792.166p 0 793.877p 0 793.878p 10000.0u 793.879p 0 802.742p 0 802.743p 10000.0u 802.744p 0 810.806p 0 810.807p 10000.0u 810.808p 0 811.151p 0 811.152p 10000.0u 811.153p 0 814.904p 0 814.905p 10000.0u 814.906p 0 825.695p 0 825.696p 10000.0u 825.697p 0 865.76p 0 865.761p 10000.0u 865.762p 0 866.054p 0 866.055p 10000.0u 866.056p 0 869.129p 0 869.13p 10000.0u 869.131p 0 870.305p 0 870.306p 10000.0u 870.307p 0 870.404p 0 870.405p 10000.0u 870.406p 0 882.791p 0 882.792p 10000.0u 882.793p 0 886.178p 0 886.179p 10000.0u 886.18p 0 888.527p 0 888.528p 10000.0u 888.529p 0 888.761p 0 888.762p 10000.0u 888.763p 0 913.322p 0 913.323p 10000.0u 913.324p 0 913.454p 0 913.455p 10000.0u 913.456p 0 955.151p 0 955.152p 10000.0u 955.153p 0 958.808p 0 958.809p 10000.0u 958.81p 0 969.278p 0 969.279p 10000.0u 969.28p 0 977.099p 0 977.1p 10000.0u 977.101p 0 978.602p 0 978.603p 10000.0u 978.604p 0)
IIN44 0 45 pwl(0 0 27.764p 0 27.765p 10000.0u 27.766p 0 34.94p 0 34.941p 10000.0u 34.942p 0 42.98p 0 42.981p 10000.0u 42.982p 0 49.937p 0 49.938p 10000.0u 49.939p 0 58.97p 0 58.971p 10000.0u 58.972p 0 76.355p 0 76.356p 10000.0u 76.357p 0 85.514p 0 85.515p 10000.0u 85.516p 0 100.499p 0 100.5p 10000.0u 100.501p 0 100.649p 0 100.65p 10000.0u 100.651p 0 116.435p 0 116.436p 10000.0u 116.437p 0 116.816p 0 116.817p 10000.0u 116.818p 0 131.024p 0 131.025p 10000.0u 131.026p 0 134.477p 0 134.478p 10000.0u 134.479p 0 142.535p 0 142.536p 10000.0u 142.537p 0 149.21p 0 149.211p 10000.0u 149.212p 0 158.075p 0 158.076p 10000.0u 158.077p 0 159.146p 0 159.147p 10000.0u 159.148p 0 167.153p 0 167.154p 10000.0u 167.155p 0 173.132p 0 173.133p 10000.0u 173.134p 0 176.066p 0 176.067p 10000.0u 176.068p 0 179.906p 0 179.907p 10000.0u 179.908p 0 188.915p 0 188.916p 10000.0u 188.917p 0 198.2p 0 198.201p 10000.0u 198.202p 0 207.971p 0 207.972p 10000.0u 207.973p 0 208.43p 0 208.431p 10000.0u 208.432p 0 217.148p 0 217.149p 10000.0u 217.15p 0 226.796p 0 226.797p 10000.0u 226.798p 0 232.439p 0 232.44p 10000.0u 232.441p 0 257.408p 0 257.409p 10000.0u 257.41p 0 257.924p 0 257.925p 10000.0u 257.926p 0 261.542p 0 261.543p 10000.0u 261.544p 0 283.571p 0 283.572p 10000.0u 283.573p 0 288.863p 0 288.864p 10000.0u 288.865p 0 304.778p 0 304.779p 10000.0u 304.78p 0 320.366p 0 320.367p 10000.0u 320.368p 0 324.89p 0 324.891p 10000.0u 324.892p 0 331.385p 0 331.386p 10000.0u 331.387p 0 349.499p 0 349.5p 10000.0u 349.501p 0 356.81p 0 356.811p 10000.0u 356.812p 0 358.52p 0 358.521p 10000.0u 358.522p 0 358.952p 0 358.953p 10000.0u 358.954p 0 369.698p 0 369.699p 10000.0u 369.7p 0 386.711p 0 386.712p 10000.0u 386.713p 0 400.952p 0 400.953p 10000.0u 400.954p 0 404.585p 0 404.586p 10000.0u 404.587p 0 413.393p 0 413.394p 10000.0u 413.395p 0 416.816p 0 416.817p 10000.0u 416.818p 0 450.41p 0 450.411p 10000.0u 450.412p 0 470.354p 0 470.355p 10000.0u 470.356p 0 472.106p 0 472.107p 10000.0u 472.108p 0 474.86p 0 474.861p 10000.0u 474.862p 0 485.201p 0 485.202p 10000.0u 485.203p 0 495.092p 0 495.093p 10000.0u 495.094p 0 504.671p 0 504.672p 10000.0u 504.673p 0 509.378p 0 509.379p 10000.0u 509.38p 0 516.254p 0 516.255p 10000.0u 516.256p 0 517.961p 0 517.962p 10000.0u 517.963p 0 533.72p 0 533.721p 10000.0u 533.722p 0 538.643p 0 538.644p 10000.0u 538.645p 0 540.515p 0 540.516p 10000.0u 540.517p 0 551.747p 0 551.748p 10000.0u 551.749p 0 573.767p 0 573.768p 10000.0u 573.769p 0 575.936p 0 575.937p 10000.0u 575.938p 0 577.292p 0 577.293p 10000.0u 577.294p 0 584.291p 0 584.292p 10000.0u 584.293p 0 588.899p 0 588.9p 10000.0u 588.901p 0 594.824p 0 594.825p 10000.0u 594.826p 0 612.452p 0 612.453p 10000.0u 612.454p 0 624.824p 0 624.825p 10000.0u 624.826p 0 636.29p 0 636.291p 10000.0u 636.292p 0 638.72p 0 638.721p 10000.0u 638.722p 0 639.239p 0 639.24p 10000.0u 639.241p 0 666.476p 0 666.477p 10000.0u 666.478p 0 669.083p 0 669.084p 10000.0u 669.085p 0 675.38p 0 675.381p 10000.0u 675.382p 0 678.206p 0 678.207p 10000.0u 678.208p 0 694.919p 0 694.92p 10000.0u 694.921p 0 715.64p 0 715.641p 10000.0u 715.642p 0 718.727p 0 718.728p 10000.0u 718.729p 0 740.096p 0 740.097p 10000.0u 740.098p 0 746.846p 0 746.847p 10000.0u 746.848p 0 771.941p 0 771.942p 10000.0u 771.943p 0 792.602p 0 792.603p 10000.0u 792.604p 0 800.153p 0 800.154p 10000.0u 800.155p 0 804.212p 0 804.213p 10000.0u 804.214p 0 805.058p 0 805.059p 10000.0u 805.06p 0 816.032p 0 816.033p 10000.0u 816.034p 0 821.969p 0 821.97p 10000.0u 821.971p 0 836.672p 0 836.673p 10000.0u 836.674p 0 838.964p 0 838.965p 10000.0u 838.966p 0 853.001p 0 853.002p 10000.0u 853.003p 0 864.836p 0 864.837p 10000.0u 864.838p 0 912.206p 0 912.207p 10000.0u 912.208p 0 931.748p 0 931.749p 10000.0u 931.75p 0 934.967p 0 934.968p 10000.0u 934.969p 0 946.643p 0 946.644p 10000.0u 946.645p 0 966.053p 0 966.054p 10000.0u 966.055p 0 975.701p 0 975.702p 10000.0u 975.703p 0 983.189p 0 983.19p 10000.0u 983.191p 0 988.181p 0 988.182p 10000.0u 988.183p 0 998.183p 0 998.184p 10000.0u 998.185p 0)
IIN45 0 46 pwl(0 0 3.617p 0 3.618p 10000.0u 3.619p 0 31.235p 0 31.236p 10000.0u 31.237p 0 63.392p 0 63.393p 10000.0u 63.394p 0 66.08p 0 66.081p 10000.0u 66.082p 0 92.375p 0 92.376p 10000.0u 92.377p 0 133.757p 0 133.758p 10000.0u 133.759p 0 142.631p 0 142.632p 10000.0u 142.633p 0 145.784p 0 145.785p 10000.0u 145.786p 0 165.659p 0 165.66p 10000.0u 165.661p 0 171.656p 0 171.657p 10000.0u 171.658p 0 173.12p 0 173.121p 10000.0u 173.122p 0 202.748p 0 202.749p 10000.0u 202.75p 0 210.713p 0 210.714p 10000.0u 210.715p 0 232.388p 0 232.389p 10000.0u 232.39p 0 251.849p 0 251.85p 10000.0u 251.851p 0 251.873p 0 251.874p 10000.0u 251.875p 0 254.135p 0 254.136p 10000.0u 254.137p 0 275.42p 0 275.421p 10000.0u 275.422p 0 275.549p 0 275.55p 10000.0u 275.551p 0 275.996p 0 275.997p 10000.0u 275.998p 0 281.414p 0 281.415p 10000.0u 281.416p 0 291.038p 0 291.039p 10000.0u 291.04p 0 294.38p 0 294.381p 10000.0u 294.382p 0 300.923p 0 300.924p 10000.0u 300.925p 0 323.438p 0 323.439p 10000.0u 323.44p 0 338.372p 0 338.373p 10000.0u 338.374p 0 344.171p 0 344.172p 10000.0u 344.173p 0 350.012p 0 350.013p 10000.0u 350.014p 0 367.106p 0 367.107p 10000.0u 367.108p 0 367.514p 0 367.515p 10000.0u 367.516p 0 377.075p 0 377.076p 10000.0u 377.077p 0 379.424p 0 379.425p 10000.0u 379.426p 0 391.175p 0 391.176p 10000.0u 391.177p 0 393.953p 0 393.954p 10000.0u 393.955p 0 395.54p 0 395.541p 10000.0u 395.542p 0 400.583p 0 400.584p 10000.0u 400.585p 0 410.258p 0 410.259p 10000.0u 410.26p 0 454.037p 0 454.038p 10000.0u 454.039p 0 467.702p 0 467.703p 10000.0u 467.704p 0 479.696p 0 479.697p 10000.0u 479.698p 0 481.226p 0 481.227p 10000.0u 481.228p 0 490.844p 0 490.845p 10000.0u 490.846p 0 491.513p 0 491.514p 10000.0u 491.515p 0 492.482p 0 492.483p 10000.0u 492.484p 0 502.628p 0 502.629p 10000.0u 502.63p 0 513.281p 0 513.282p 10000.0u 513.283p 0 533.06p 0 533.061p 10000.0u 533.062p 0 558.185p 0 558.186p 10000.0u 558.187p 0 568.151p 0 568.152p 10000.0u 568.153p 0 568.622p 0 568.623p 10000.0u 568.624p 0 574.901p 0 574.902p 10000.0u 574.903p 0 579.452p 0 579.453p 10000.0u 579.454p 0 586.616p 0 586.617p 10000.0u 586.618p 0 607.55p 0 607.551p 10000.0u 607.552p 0 615.812p 0 615.813p 10000.0u 615.814p 0 622.979p 0 622.98p 10000.0u 622.981p 0 631.979p 0 631.98p 10000.0u 631.981p 0 644.828p 0 644.829p 10000.0u 644.83p 0 667.256p 0 667.257p 10000.0u 667.258p 0 668.06p 0 668.061p 10000.0u 668.062p 0 672.536p 0 672.537p 10000.0u 672.538p 0 679.814p 0 679.815p 10000.0u 679.816p 0 691.094p 0 691.095p 10000.0u 691.096p 0 698.669p 0 698.67p 10000.0u 698.671p 0 702.671p 0 702.672p 10000.0u 702.673p 0 711.605p 0 711.606p 10000.0u 711.607p 0 726.845p 0 726.846p 10000.0u 726.847p 0 749.708p 0 749.709p 10000.0u 749.71p 0 772.166p 0 772.167p 10000.0u 772.168p 0 777.311p 0 777.312p 10000.0u 777.313p 0 783.092p 0 783.093p 10000.0u 783.094p 0 800.327p 0 800.328p 10000.0u 800.329p 0 800.78p 0 800.781p 10000.0u 800.782p 0 803.516p 0 803.517p 10000.0u 803.518p 0 816.374p 0 816.375p 10000.0u 816.376p 0 817.448p 0 817.449p 10000.0u 817.45p 0 820.004p 0 820.005p 10000.0u 820.006p 0 835.943p 0 835.944p 10000.0u 835.945p 0 836.675p 0 836.676p 10000.0u 836.677p 0 854.159p 0 854.16p 10000.0u 854.161p 0 854.306p 0 854.307p 10000.0u 854.308p 0 863.441p 0 863.442p 10000.0u 863.443p 0 863.567p 0 863.568p 10000.0u 863.569p 0 870.791p 0 870.792p 10000.0u 870.793p 0 871.832p 0 871.833p 10000.0u 871.834p 0 882.602p 0 882.603p 10000.0u 882.604p 0 883.853p 0 883.854p 10000.0u 883.855p 0 889.298p 0 889.299p 10000.0u 889.3p 0 895.076p 0 895.077p 10000.0u 895.078p 0 895.391p 0 895.392p 10000.0u 895.393p 0 898.82p 0 898.821p 10000.0u 898.822p 0 901.73p 0 901.731p 10000.0u 901.732p 0 902.357p 0 902.358p 10000.0u 902.359p 0 903.029p 0 903.03p 10000.0u 903.031p 0 904.64p 0 904.641p 10000.0u 904.642p 0 922.097p 0 922.098p 10000.0u 922.099p 0 933.485p 0 933.486p 10000.0u 933.487p 0 934.025p 0 934.026p 10000.0u 934.027p 0 938.027p 0 938.028p 10000.0u 938.029p 0 938.444p 0 938.445p 10000.0u 938.446p 0 957.905p 0 957.906p 10000.0u 957.907p 0)
IIN46 0 47 pwl(0 0 21.002p 0 21.003p 10000.0u 21.004p 0 37.892p 0 37.893p 10000.0u 37.894p 0 42.545p 0 42.546p 10000.0u 42.547p 0 47.228p 0 47.229p 10000.0u 47.23p 0 52.073p 0 52.074p 10000.0u 52.075p 0 56.534p 0 56.535p 10000.0u 56.536p 0 57.83p 0 57.831p 10000.0u 57.832p 0 58.445p 0 58.446p 10000.0u 58.447p 0 58.67p 0 58.671p 10000.0u 58.672p 0 68.375p 0 68.376p 10000.0u 68.377p 0 80.852p 0 80.853p 10000.0u 80.854p 0 84.242p 0 84.243p 10000.0u 84.244p 0 88.172p 0 88.173p 10000.0u 88.174p 0 88.205p 0 88.206p 10000.0u 88.207p 0 90.602p 0 90.603p 10000.0u 90.604p 0 93.902p 0 93.903p 10000.0u 93.904p 0 99.98p 0 99.981p 10000.0u 99.982p 0 109.181p 0 109.182p 10000.0u 109.183p 0 113.684p 0 113.685p 10000.0u 113.686p 0 119.078p 0 119.079p 10000.0u 119.08p 0 137.825p 0 137.826p 10000.0u 137.827p 0 142.037p 0 142.038p 10000.0u 142.039p 0 157.976p 0 157.977p 10000.0u 157.978p 0 174.155p 0 174.156p 10000.0u 174.157p 0 176.294p 0 176.295p 10000.0u 176.296p 0 186.527p 0 186.528p 10000.0u 186.529p 0 194.576p 0 194.577p 10000.0u 194.578p 0 203.681p 0 203.682p 10000.0u 203.683p 0 212.159p 0 212.16p 10000.0u 212.161p 0 227.615p 0 227.616p 10000.0u 227.617p 0 241.457p 0 241.458p 10000.0u 241.459p 0 244.907p 0 244.908p 10000.0u 244.909p 0 245.882p 0 245.883p 10000.0u 245.884p 0 247.76p 0 247.761p 10000.0u 247.762p 0 249.92p 0 249.921p 10000.0u 249.922p 0 260.48p 0 260.481p 10000.0u 260.482p 0 268.376p 0 268.377p 10000.0u 268.378p 0 271.775p 0 271.776p 10000.0u 271.777p 0 283.712p 0 283.713p 10000.0u 283.714p 0 290.342p 0 290.343p 10000.0u 290.344p 0 298.715p 0 298.716p 10000.0u 298.717p 0 313.994p 0 313.995p 10000.0u 313.996p 0 329.921p 0 329.922p 10000.0u 329.923p 0 342.965p 0 342.966p 10000.0u 342.967p 0 355.817p 0 355.818p 10000.0u 355.819p 0 363.518p 0 363.519p 10000.0u 363.52p 0 388.058p 0 388.059p 10000.0u 388.06p 0 388.853p 0 388.854p 10000.0u 388.855p 0 397.187p 0 397.188p 10000.0u 397.189p 0 402.224p 0 402.225p 10000.0u 402.226p 0 404.78p 0 404.781p 10000.0u 404.782p 0 419.804p 0 419.805p 10000.0u 419.806p 0 433.622p 0 433.623p 10000.0u 433.624p 0 437.318p 0 437.319p 10000.0u 437.32p 0 452.924p 0 452.925p 10000.0u 452.926p 0 454.91p 0 454.911p 10000.0u 454.912p 0 468.632p 0 468.633p 10000.0u 468.634p 0 470.429p 0 470.43p 10000.0u 470.431p 0 488.978p 0 488.979p 10000.0u 488.98p 0 490.169p 0 490.17p 10000.0u 490.171p 0 499.607p 0 499.608p 10000.0u 499.609p 0 500.867p 0 500.868p 10000.0u 500.869p 0 506.861p 0 506.862p 10000.0u 506.863p 0 511.016p 0 511.017p 10000.0u 511.018p 0 523.694p 0 523.695p 10000.0u 523.696p 0 544.511p 0 544.512p 10000.0u 544.513p 0 556.505p 0 556.506p 10000.0u 556.507p 0 569.126p 0 569.127p 10000.0u 569.128p 0 591.38p 0 591.381p 10000.0u 591.382p 0 598.652p 0 598.653p 10000.0u 598.654p 0 599.705p 0 599.706p 10000.0u 599.707p 0 620.132p 0 620.133p 10000.0u 620.134p 0 641.528p 0 641.529p 10000.0u 641.53p 0 648.29p 0 648.291p 10000.0u 648.292p 0 667.205p 0 667.206p 10000.0u 667.207p 0 674.393p 0 674.394p 10000.0u 674.395p 0 685.16p 0 685.161p 10000.0u 685.162p 0 689.309p 0 689.31p 10000.0u 689.311p 0 732.611p 0 732.612p 10000.0u 732.613p 0 741.455p 0 741.456p 10000.0u 741.457p 0 741.632p 0 741.633p 10000.0u 741.634p 0 755.846p 0 755.847p 10000.0u 755.848p 0 763.487p 0 763.488p 10000.0u 763.489p 0 768.926p 0 768.927p 10000.0u 768.928p 0 770.357p 0 770.358p 10000.0u 770.359p 0 771.329p 0 771.33p 10000.0u 771.331p 0 772.013p 0 772.014p 10000.0u 772.015p 0 776.981p 0 776.982p 10000.0u 776.983p 0 786.209p 0 786.21p 10000.0u 786.211p 0 808.331p 0 808.332p 10000.0u 808.333p 0 816.92p 0 816.921p 10000.0u 816.922p 0 826.637p 0 826.638p 10000.0u 826.639p 0 837.407p 0 837.408p 10000.0u 837.409p 0 844.925p 0 844.926p 10000.0u 844.927p 0 846.707p 0 846.708p 10000.0u 846.709p 0 850.439p 0 850.44p 10000.0u 850.441p 0 852.824p 0 852.825p 10000.0u 852.826p 0 891.863p 0 891.864p 10000.0u 891.865p 0 895.007p 0 895.008p 10000.0u 895.009p 0 898.232p 0 898.233p 10000.0u 898.234p 0 919.268p 0 919.269p 10000.0u 919.27p 0 927.695p 0 927.696p 10000.0u 927.697p 0 958.331p 0 958.332p 10000.0u 958.333p 0 987.023p 0 987.024p 10000.0u 987.025p 0 992.579p 0 992.58p 10000.0u 992.581p 0 993.41p 0 993.411p 10000.0u 993.412p 0 999.2p 0 999.201p 10000.0u 999.202p 0)
IIN47 0 48 pwl(0 0 16.22p 0 16.221p 10000.0u 16.222p 0 26.519p 0 26.52p 10000.0u 26.521p 0 31.424p 0 31.425p 10000.0u 31.426p 0 31.898p 0 31.899p 10000.0u 31.9p 0 43.934p 0 43.935p 10000.0u 43.936p 0 52.415p 0 52.416p 10000.0u 52.417p 0 76.616p 0 76.617p 10000.0u 76.618p 0 95.744p 0 95.745p 10000.0u 95.746p 0 101.888p 0 101.889p 10000.0u 101.89p 0 129.341p 0 129.342p 10000.0u 129.343p 0 130.367p 0 130.368p 10000.0u 130.369p 0 138.224p 0 138.225p 10000.0u 138.226p 0 152.252p 0 152.253p 10000.0u 152.254p 0 163.25p 0 163.251p 10000.0u 163.252p 0 171.464p 0 171.465p 10000.0u 171.466p 0 178.283p 0 178.284p 10000.0u 178.285p 0 199.961p 0 199.962p 10000.0u 199.963p 0 201.605p 0 201.606p 10000.0u 201.607p 0 205.949p 0 205.95p 10000.0u 205.951p 0 234.656p 0 234.657p 10000.0u 234.658p 0 238.112p 0 238.113p 10000.0u 238.114p 0 239.102p 0 239.103p 10000.0u 239.104p 0 279.221p 0 279.222p 10000.0u 279.223p 0 295.727p 0 295.728p 10000.0u 295.729p 0 322.088p 0 322.089p 10000.0u 322.09p 0 323.108p 0 323.109p 10000.0u 323.11p 0 323.81p 0 323.811p 10000.0u 323.812p 0 328.922p 0 328.923p 10000.0u 328.924p 0 329.072p 0 329.073p 10000.0u 329.074p 0 337.847p 0 337.848p 10000.0u 337.849p 0 338.945p 0 338.946p 10000.0u 338.947p 0 347.522p 0 347.523p 10000.0u 347.524p 0 360.866p 0 360.867p 10000.0u 360.868p 0 362.432p 0 362.433p 10000.0u 362.434p 0 380.576p 0 380.577p 10000.0u 380.578p 0 385.433p 0 385.434p 10000.0u 385.435p 0 385.763p 0 385.764p 10000.0u 385.765p 0 404.54p 0 404.541p 10000.0u 404.542p 0 412.508p 0 412.509p 10000.0u 412.51p 0 423.038p 0 423.039p 10000.0u 423.04p 0 438.155p 0 438.156p 10000.0u 438.157p 0 439.475p 0 439.476p 10000.0u 439.477p 0 441.71p 0 441.711p 10000.0u 441.712p 0 453.716p 0 453.717p 10000.0u 453.718p 0 464.345p 0 464.346p 10000.0u 464.347p 0 472.382p 0 472.383p 10000.0u 472.384p 0 482.63p 0 482.631p 10000.0u 482.632p 0 487.877p 0 487.878p 10000.0u 487.879p 0 499.718p 0 499.719p 10000.0u 499.72p 0 501.545p 0 501.546p 10000.0u 501.547p 0 517.379p 0 517.38p 10000.0u 517.381p 0 520.595p 0 520.596p 10000.0u 520.597p 0 537.038p 0 537.039p 10000.0u 537.04p 0 549.263p 0 549.264p 10000.0u 549.265p 0 549.596p 0 549.597p 10000.0u 549.598p 0 553.229p 0 553.23p 10000.0u 553.231p 0 567.884p 0 567.885p 10000.0u 567.886p 0 575.918p 0 575.919p 10000.0u 575.92p 0 578.957p 0 578.958p 10000.0u 578.959p 0 587.213p 0 587.214p 10000.0u 587.215p 0 623.924p 0 623.925p 10000.0u 623.926p 0 625.166p 0 625.167p 10000.0u 625.168p 0 626.009p 0 626.01p 10000.0u 626.011p 0 634.298p 0 634.299p 10000.0u 634.3p 0 640.103p 0 640.104p 10000.0u 640.105p 0 640.106p 0 640.107p 10000.0u 640.108p 0 644.801p 0 644.802p 10000.0u 644.803p 0 646.67p 0 646.671p 10000.0u 646.672p 0 650.906p 0 650.907p 10000.0u 650.908p 0 655.016p 0 655.017p 10000.0u 655.018p 0 663.272p 0 663.273p 10000.0u 663.274p 0 664.676p 0 664.677p 10000.0u 664.678p 0 665.813p 0 665.814p 10000.0u 665.815p 0 667.439p 0 667.44p 10000.0u 667.441p 0 674.816p 0 674.817p 10000.0u 674.818p 0 689.117p 0 689.118p 10000.0u 689.119p 0 704.036p 0 704.037p 10000.0u 704.038p 0 708.056p 0 708.057p 10000.0u 708.058p 0 711.26p 0 711.261p 10000.0u 711.262p 0 715.151p 0 715.152p 10000.0u 715.153p 0 744.911p 0 744.912p 10000.0u 744.913p 0 761.669p 0 761.67p 10000.0u 761.671p 0 766.193p 0 766.194p 10000.0u 766.195p 0 769.448p 0 769.449p 10000.0u 769.45p 0 771.734p 0 771.735p 10000.0u 771.736p 0 775.322p 0 775.323p 10000.0u 775.324p 0 803.942p 0 803.943p 10000.0u 803.944p 0 813.341p 0 813.342p 10000.0u 813.343p 0 840.071p 0 840.072p 10000.0u 840.073p 0 855.857p 0 855.858p 10000.0u 855.859p 0 867.911p 0 867.912p 10000.0u 867.913p 0 878.399p 0 878.4p 10000.0u 878.401p 0 886.565p 0 886.566p 10000.0u 886.567p 0 898.106p 0 898.107p 10000.0u 898.108p 0 904.139p 0 904.14p 10000.0u 904.141p 0 906.545p 0 906.546p 10000.0u 906.547p 0 927.338p 0 927.339p 10000.0u 927.34p 0 950.942p 0 950.943p 10000.0u 950.944p 0 969.278p 0 969.279p 10000.0u 969.28p 0 978.908p 0 978.909p 10000.0u 978.91p 0 979.406p 0 979.407p 10000.0u 979.408p 0 983.018p 0 983.019p 10000.0u 983.02p 0 984.032p 0 984.033p 10000.0u 984.034p 0 992.204p 0 992.205p 10000.0u 992.206p 0)
IIN48 0 49 pwl(0 0 4.658p 0 4.659p 10000.0u 4.66p 0 5.561p 0 5.562p 10000.0u 5.563p 0 18.191p 0 18.192p 10000.0u 18.193p 0 21.881p 0 21.882p 10000.0u 21.883p 0 24.581p 0 24.582p 10000.0u 24.583p 0 25.256p 0 25.257p 10000.0u 25.258p 0 27.086p 0 27.087p 10000.0u 27.088p 0 65.66p 0 65.661p 10000.0u 65.662p 0 75.272p 0 75.273p 10000.0u 75.274p 0 80.897p 0 80.898p 10000.0u 80.899p 0 96.788p 0 96.789p 10000.0u 96.79p 0 99.821p 0 99.822p 10000.0u 99.823p 0 113.474p 0 113.475p 10000.0u 113.476p 0 119.129p 0 119.13p 10000.0u 119.131p 0 140.225p 0 140.226p 10000.0u 140.227p 0 150.53p 0 150.531p 10000.0u 150.532p 0 164.096p 0 164.097p 10000.0u 164.098p 0 178.667p 0 178.668p 10000.0u 178.669p 0 180.806p 0 180.807p 10000.0u 180.808p 0 188.258p 0 188.259p 10000.0u 188.26p 0 216.734p 0 216.735p 10000.0u 216.736p 0 220.508p 0 220.509p 10000.0u 220.51p 0 226.295p 0 226.296p 10000.0u 226.297p 0 227.885p 0 227.886p 10000.0u 227.887p 0 266.504p 0 266.505p 10000.0u 266.506p 0 273.797p 0 273.798p 10000.0u 273.799p 0 282.494p 0 282.495p 10000.0u 282.496p 0 283.805p 0 283.806p 10000.0u 283.807p 0 284.216p 0 284.217p 10000.0u 284.218p 0 284.726p 0 284.727p 10000.0u 284.728p 0 288.173p 0 288.174p 10000.0u 288.175p 0 294.581p 0 294.582p 10000.0u 294.583p 0 298.106p 0 298.107p 10000.0u 298.108p 0 307.616p 0 307.617p 10000.0u 307.618p 0 316.115p 0 316.116p 10000.0u 316.117p 0 325.388p 0 325.389p 10000.0u 325.39p 0 338.558p 0 338.559p 10000.0u 338.56p 0 345.716p 0 345.717p 10000.0u 345.718p 0 387.059p 0 387.06p 10000.0u 387.061p 0 432.428p 0 432.429p 10000.0u 432.43p 0 439.277p 0 439.278p 10000.0u 439.279p 0 449.588p 0 449.589p 10000.0u 449.59p 0 449.963p 0 449.964p 10000.0u 449.965p 0 460.295p 0 460.296p 10000.0u 460.297p 0 469.301p 0 469.302p 10000.0u 469.303p 0 470.198p 0 470.199p 10000.0u 470.2p 0 477.8p 0 477.801p 10000.0u 477.802p 0 493.64p 0 493.641p 10000.0u 493.642p 0 496.856p 0 496.857p 10000.0u 496.858p 0 499.382p 0 499.383p 10000.0u 499.384p 0 502.376p 0 502.377p 10000.0u 502.378p 0 507.626p 0 507.627p 10000.0u 507.628p 0 520.061p 0 520.062p 10000.0u 520.063p 0 520.901p 0 520.902p 10000.0u 520.903p 0 528.92p 0 528.921p 10000.0u 528.922p 0 566.735p 0 566.736p 10000.0u 566.737p 0 568.853p 0 568.854p 10000.0u 568.855p 0 569.702p 0 569.703p 10000.0u 569.704p 0 574.895p 0 574.896p 10000.0u 574.897p 0 596.945p 0 596.946p 10000.0u 596.947p 0 610.217p 0 610.218p 10000.0u 610.219p 0 635.558p 0 635.559p 10000.0u 635.56p 0 638.462p 0 638.463p 10000.0u 638.464p 0 640.655p 0 640.656p 10000.0u 640.657p 0 654.83p 0 654.831p 10000.0u 654.832p 0 667.079p 0 667.08p 10000.0u 667.081p 0 682.271p 0 682.272p 10000.0u 682.273p 0 691.487p 0 691.488p 10000.0u 691.489p 0 693.56p 0 693.561p 10000.0u 693.562p 0 704.921p 0 704.922p 10000.0u 704.923p 0 713.447p 0 713.448p 10000.0u 713.449p 0 723.68p 0 723.681p 10000.0u 723.682p 0 735.5p 0 735.501p 10000.0u 735.502p 0 736.304p 0 736.305p 10000.0u 736.306p 0 752.36p 0 752.361p 10000.0u 752.362p 0 763.412p 0 763.413p 10000.0u 763.414p 0 782.585p 0 782.586p 10000.0u 782.587p 0 789.509p 0 789.51p 10000.0u 789.511p 0 800.642p 0 800.643p 10000.0u 800.644p 0 801.701p 0 801.702p 10000.0u 801.703p 0 811.664p 0 811.665p 10000.0u 811.666p 0 813.908p 0 813.909p 10000.0u 813.91p 0 856.379p 0 856.38p 10000.0u 856.381p 0 885.194p 0 885.195p 10000.0u 885.196p 0 887.618p 0 887.619p 10000.0u 887.62p 0 889.625p 0 889.626p 10000.0u 889.627p 0 890.822p 0 890.823p 10000.0u 890.824p 0 892.694p 0 892.695p 10000.0u 892.696p 0 893.69p 0 893.691p 10000.0u 893.692p 0 901.466p 0 901.467p 10000.0u 901.468p 0 910.742p 0 910.743p 10000.0u 910.744p 0 911.999p 0 912.0p 10000.0u 912.001p 0 913.982p 0 913.983p 10000.0u 913.984p 0 949.085p 0 949.086p 10000.0u 949.087p 0 950.135p 0 950.136p 10000.0u 950.137p 0 955.796p 0 955.797p 10000.0u 955.798p 0 970.721p 0 970.722p 10000.0u 970.723p 0 977.474p 0 977.475p 10000.0u 977.476p 0 983.348p 0 983.349p 10000.0u 983.35p 0 988.235p 0 988.236p 10000.0u 988.237p 0 989.198p 0 989.199p 10000.0u 989.2p 0)
IIN49 0 50 pwl(0 0 37.511p 0 37.512p 10000.0u 37.513p 0 49.73p 0 49.731p 10000.0u 49.732p 0 50.861p 0 50.862p 10000.0u 50.863p 0 54.602p 0 54.603p 10000.0u 54.604p 0 55.214p 0 55.215p 10000.0u 55.216p 0 59.192p 0 59.193p 10000.0u 59.194p 0 84.5p 0 84.501p 10000.0u 84.502p 0 89.414p 0 89.415p 10000.0u 89.416p 0 92.045p 0 92.046p 10000.0u 92.047p 0 93.857p 0 93.858p 10000.0u 93.859p 0 94.217p 0 94.218p 10000.0u 94.219p 0 105.254p 0 105.255p 10000.0u 105.256p 0 110.915p 0 110.916p 10000.0u 110.917p 0 113.249p 0 113.25p 10000.0u 113.251p 0 117.875p 0 117.876p 10000.0u 117.877p 0 140.909p 0 140.91p 10000.0u 140.911p 0 146.924p 0 146.925p 10000.0u 146.926p 0 149.567p 0 149.568p 10000.0u 149.569p 0 156.518p 0 156.519p 10000.0u 156.52p 0 181.274p 0 181.275p 10000.0u 181.276p 0 192.8p 0 192.801p 10000.0u 192.802p 0 192.848p 0 192.849p 10000.0u 192.85p 0 197.714p 0 197.715p 10000.0u 197.716p 0 200.732p 0 200.733p 10000.0u 200.734p 0 215.699p 0 215.7p 10000.0u 215.701p 0 215.987p 0 215.988p 10000.0u 215.989p 0 245.489p 0 245.49p 10000.0u 245.491p 0 246.539p 0 246.54p 10000.0u 246.541p 0 267.149p 0 267.15p 10000.0u 267.151p 0 284.675p 0 284.676p 10000.0u 284.677p 0 299.882p 0 299.883p 10000.0u 299.884p 0 301.592p 0 301.593p 10000.0u 301.594p 0 307.697p 0 307.698p 10000.0u 307.699p 0 311.876p 0 311.877p 10000.0u 311.878p 0 326.609p 0 326.61p 10000.0u 326.611p 0 342.563p 0 342.564p 10000.0u 342.565p 0 343.16p 0 343.161p 10000.0u 343.162p 0 346.841p 0 346.842p 10000.0u 346.843p 0 383.375p 0 383.376p 10000.0u 383.377p 0 385.514p 0 385.515p 10000.0u 385.516p 0 400.376p 0 400.377p 10000.0u 400.378p 0 401.327p 0 401.328p 10000.0u 401.329p 0 402.53p 0 402.531p 10000.0u 402.532p 0 426.023p 0 426.024p 10000.0u 426.025p 0 439.097p 0 439.098p 10000.0u 439.099p 0 439.406p 0 439.407p 10000.0u 439.408p 0 442.808p 0 442.809p 10000.0u 442.81p 0 453.62p 0 453.621p 10000.0u 453.622p 0 463.565p 0 463.566p 10000.0u 463.567p 0 465.845p 0 465.846p 10000.0u 465.847p 0 467.177p 0 467.178p 10000.0u 467.179p 0 482.147p 0 482.148p 10000.0u 482.149p 0 497.492p 0 497.493p 10000.0u 497.494p 0 500.978p 0 500.979p 10000.0u 500.98p 0 507.98p 0 507.981p 10000.0u 507.982p 0 509.936p 0 509.937p 10000.0u 509.938p 0 526.37p 0 526.371p 10000.0u 526.372p 0 527.243p 0 527.244p 10000.0u 527.245p 0 536.744p 0 536.745p 10000.0u 536.746p 0 542.522p 0 542.523p 10000.0u 542.524p 0 547.337p 0 547.338p 10000.0u 547.339p 0 552.725p 0 552.726p 10000.0u 552.727p 0 560.81p 0 560.811p 10000.0u 560.812p 0 561.71p 0 561.711p 10000.0u 561.712p 0 571.19p 0 571.191p 10000.0u 571.192p 0 587.219p 0 587.22p 10000.0u 587.221p 0 592.208p 0 592.209p 10000.0u 592.21p 0 599.552p 0 599.553p 10000.0u 599.554p 0 608.153p 0 608.154p 10000.0u 608.155p 0 609.08p 0 609.081p 10000.0u 609.082p 0 617.36p 0 617.361p 10000.0u 617.362p 0 629.579p 0 629.58p 10000.0u 629.581p 0 630.14p 0 630.141p 10000.0u 630.142p 0 632.57p 0 632.571p 10000.0u 632.572p 0 638.024p 0 638.025p 10000.0u 638.026p 0 648.221p 0 648.222p 10000.0u 648.223p 0 658.391p 0 658.392p 10000.0u 658.393p 0 658.958p 0 658.959p 10000.0u 658.96p 0 665.963p 0 665.964p 10000.0u 665.965p 0 667.793p 0 667.794p 10000.0u 667.795p 0 677.348p 0 677.349p 10000.0u 677.35p 0 691.001p 0 691.002p 10000.0u 691.003p 0 719.867p 0 719.868p 10000.0u 719.869p 0 720.773p 0 720.774p 10000.0u 720.775p 0 724.133p 0 724.134p 10000.0u 724.135p 0 735.407p 0 735.408p 10000.0u 735.409p 0 748.217p 0 748.218p 10000.0u 748.219p 0 750.065p 0 750.066p 10000.0u 750.067p 0 761.486p 0 761.487p 10000.0u 761.488p 0 762.356p 0 762.357p 10000.0u 762.358p 0 764.141p 0 764.142p 10000.0u 764.143p 0 765.197p 0 765.198p 10000.0u 765.199p 0 772.934p 0 772.935p 10000.0u 772.936p 0 774.995p 0 774.996p 10000.0u 774.997p 0 781.289p 0 781.29p 10000.0u 781.291p 0 782.39p 0 782.391p 10000.0u 782.392p 0 789.608p 0 789.609p 10000.0u 789.61p 0 793.103p 0 793.104p 10000.0u 793.105p 0 803.693p 0 803.694p 10000.0u 803.695p 0 807.227p 0 807.228p 10000.0u 807.229p 0 824.681p 0 824.682p 10000.0u 824.683p 0 840.473p 0 840.474p 10000.0u 840.475p 0 840.623p 0 840.624p 10000.0u 840.625p 0 850.472p 0 850.473p 10000.0u 850.474p 0 851.624p 0 851.625p 10000.0u 851.626p 0 867.416p 0 867.417p 10000.0u 867.418p 0 868.691p 0 868.692p 10000.0u 868.693p 0 894.137p 0 894.138p 10000.0u 894.139p 0 898.043p 0 898.044p 10000.0u 898.045p 0 900.995p 0 900.996p 10000.0u 900.997p 0 906.077p 0 906.078p 10000.0u 906.079p 0 908.546p 0 908.547p 10000.0u 908.548p 0 919.847p 0 919.848p 10000.0u 919.849p 0 930.05p 0 930.051p 10000.0u 930.052p 0 930.104p 0 930.105p 10000.0u 930.106p 0 954.134p 0 954.135p 10000.0u 954.136p 0 958.124p 0 958.125p 10000.0u 958.126p 0 974.45p 0 974.451p 10000.0u 974.452p 0 984.122p 0 984.123p 10000.0u 984.124p 0 999.437p 0 999.438p 10000.0u 999.439p 0)
IIN50 0 51 pwl(0 0 42.713p 0 42.714p 10000.0u 42.715p 0 43.892p 0 43.893p 10000.0u 43.894p 0 49.136p 0 49.137p 10000.0u 49.138p 0 52.961p 0 52.962p 10000.0u 52.963p 0 58.853p 0 58.854p 10000.0u 58.855p 0 62.669p 0 62.67p 10000.0u 62.671p 0 68.729p 0 68.73p 10000.0u 68.731p 0 71.399p 0 71.4p 10000.0u 71.401p 0 71.708p 0 71.709p 10000.0u 71.71p 0 75.209p 0 75.21p 10000.0u 75.211p 0 78.998p 0 78.999p 10000.0u 79.0p 0 104.798p 0 104.799p 10000.0u 104.8p 0 108.782p 0 108.783p 10000.0u 108.784p 0 128.777p 0 128.778p 10000.0u 128.779p 0 133.778p 0 133.779p 10000.0u 133.78p 0 136.889p 0 136.89p 10000.0u 136.891p 0 147.062p 0 147.063p 10000.0u 147.064p 0 151.181p 0 151.182p 10000.0u 151.183p 0 160.757p 0 160.758p 10000.0u 160.759p 0 172.499p 0 172.5p 10000.0u 172.501p 0 193.073p 0 193.074p 10000.0u 193.075p 0 209.348p 0 209.349p 10000.0u 209.35p 0 210.107p 0 210.108p 10000.0u 210.109p 0 212.408p 0 212.409p 10000.0u 212.41p 0 220.391p 0 220.392p 10000.0u 220.393p 0 220.55p 0 220.551p 10000.0u 220.552p 0 257.591p 0 257.592p 10000.0u 257.593p 0 259.334p 0 259.335p 10000.0u 259.336p 0 259.826p 0 259.827p 10000.0u 259.828p 0 260.006p 0 260.007p 10000.0u 260.008p 0 264.656p 0 264.657p 10000.0u 264.658p 0 268.496p 0 268.497p 10000.0u 268.498p 0 293.108p 0 293.109p 10000.0u 293.11p 0 293.744p 0 293.745p 10000.0u 293.746p 0 294.974p 0 294.975p 10000.0u 294.976p 0 308.141p 0 308.142p 10000.0u 308.143p 0 312.248p 0 312.249p 10000.0u 312.25p 0 317.864p 0 317.865p 10000.0u 317.866p 0 330.032p 0 330.033p 10000.0u 330.034p 0 344.222p 0 344.223p 10000.0u 344.224p 0 367.247p 0 367.248p 10000.0u 367.249p 0 378.11p 0 378.111p 10000.0u 378.112p 0 393.356p 0 393.357p 10000.0u 393.358p 0 395.438p 0 395.439p 10000.0u 395.44p 0 402.746p 0 402.747p 10000.0u 402.748p 0 408.041p 0 408.042p 10000.0u 408.043p 0 409.136p 0 409.137p 10000.0u 409.138p 0 414.497p 0 414.498p 10000.0u 414.499p 0 433.055p 0 433.056p 10000.0u 433.057p 0 439.652p 0 439.653p 10000.0u 439.654p 0 450.8p 0 450.801p 10000.0u 450.802p 0 455.603p 0 455.604p 10000.0u 455.605p 0 477.515p 0 477.516p 10000.0u 477.517p 0 492.65p 0 492.651p 10000.0u 492.652p 0 497.243p 0 497.244p 10000.0u 497.245p 0 498.569p 0 498.57p 10000.0u 498.571p 0 499.736p 0 499.737p 10000.0u 499.738p 0 508.1p 0 508.101p 10000.0u 508.102p 0 532.913p 0 532.914p 10000.0u 532.915p 0 551.534p 0 551.535p 10000.0u 551.536p 0 554.777p 0 554.778p 10000.0u 554.779p 0 560.363p 0 560.364p 10000.0u 560.365p 0 560.603p 0 560.604p 10000.0u 560.605p 0 574.664p 0 574.665p 10000.0u 574.666p 0 592.484p 0 592.485p 10000.0u 592.486p 0 606.329p 0 606.33p 10000.0u 606.331p 0 607.157p 0 607.158p 10000.0u 607.159p 0 607.298p 0 607.299p 10000.0u 607.3p 0 625.208p 0 625.209p 10000.0u 625.21p 0 627.413p 0 627.414p 10000.0u 627.415p 0 646.448p 0 646.449p 10000.0u 646.45p 0 650.921p 0 650.922p 10000.0u 650.923p 0 659.768p 0 659.769p 10000.0u 659.77p 0 663.452p 0 663.453p 10000.0u 663.454p 0 669.344p 0 669.345p 10000.0u 669.346p 0 679.454p 0 679.455p 10000.0u 679.456p 0 687.47p 0 687.471p 10000.0u 687.472p 0 694.322p 0 694.323p 10000.0u 694.324p 0 722.588p 0 722.589p 10000.0u 722.59p 0 724.757p 0 724.758p 10000.0u 724.759p 0 745.826p 0 745.827p 10000.0u 745.828p 0 757.259p 0 757.26p 10000.0u 757.261p 0 763.433p 0 763.434p 10000.0u 763.435p 0 776.702p 0 776.703p 10000.0u 776.704p 0 808.223p 0 808.224p 10000.0u 808.225p 0 809.999p 0 810.0p 10000.0u 810.001p 0 810.23p 0 810.231p 10000.0u 810.232p 0 823.814p 0 823.815p 10000.0u 823.816p 0 827.495p 0 827.496p 10000.0u 827.497p 0 835.277p 0 835.278p 10000.0u 835.279p 0 840.59p 0 840.591p 10000.0u 840.592p 0 849.296p 0 849.297p 10000.0u 849.298p 0 855.038p 0 855.039p 10000.0u 855.04p 0 865.367p 0 865.368p 10000.0u 865.369p 0 867.839p 0 867.84p 10000.0u 867.841p 0 878.813p 0 878.814p 10000.0u 878.815p 0 894.998p 0 894.999p 10000.0u 895.0p 0 901.7p 0 901.701p 10000.0u 901.702p 0 904.751p 0 904.752p 10000.0u 904.753p 0 921.257p 0 921.258p 10000.0u 921.259p 0 924.149p 0 924.15p 10000.0u 924.151p 0 927.791p 0 927.792p 10000.0u 927.793p 0 950.21p 0 950.211p 10000.0u 950.212p 0 956.339p 0 956.34p 10000.0u 956.341p 0 956.666p 0 956.667p 10000.0u 956.668p 0 970.379p 0 970.38p 10000.0u 970.381p 0 982.46p 0 982.461p 10000.0u 982.462p 0 994.496p 0 994.497p 10000.0u 994.498p 0)
IIN51 0 52 pwl(0 0 4.799p 0 4.8p 10000.0u 4.801p 0 12.689p 0 12.69p 10000.0u 12.691p 0 12.719p 0 12.72p 10000.0u 12.721p 0 20.771p 0 20.772p 10000.0u 20.773p 0 23.609p 0 23.61p 10000.0u 23.611p 0 27.155p 0 27.156p 10000.0u 27.157p 0 35.159p 0 35.16p 10000.0u 35.161p 0 42.566p 0 42.567p 10000.0u 42.568p 0 45.476p 0 45.477p 10000.0u 45.478p 0 51.959p 0 51.96p 10000.0u 51.961p 0 68.885p 0 68.886p 10000.0u 68.887p 0 76.172p 0 76.173p 10000.0u 76.174p 0 81.593p 0 81.594p 10000.0u 81.595p 0 90.254p 0 90.255p 10000.0u 90.256p 0 94.913p 0 94.914p 10000.0u 94.915p 0 138.68p 0 138.681p 10000.0u 138.682p 0 140.261p 0 140.262p 10000.0u 140.263p 0 153.047p 0 153.048p 10000.0u 153.049p 0 156.59p 0 156.591p 10000.0u 156.592p 0 175.598p 0 175.599p 10000.0u 175.6p 0 190.298p 0 190.299p 10000.0u 190.3p 0 191.009p 0 191.01p 10000.0u 191.011p 0 196.334p 0 196.335p 10000.0u 196.336p 0 198.812p 0 198.813p 10000.0u 198.814p 0 202.544p 0 202.545p 10000.0u 202.546p 0 204.149p 0 204.15p 10000.0u 204.151p 0 204.893p 0 204.894p 10000.0u 204.895p 0 205.289p 0 205.29p 10000.0u 205.291p 0 208.913p 0 208.914p 10000.0u 208.915p 0 212.981p 0 212.982p 10000.0u 212.983p 0 213.224p 0 213.225p 10000.0u 213.226p 0 226.925p 0 226.926p 10000.0u 226.927p 0 229.799p 0 229.8p 10000.0u 229.801p 0 265.79p 0 265.791p 10000.0u 265.792p 0 270.407p 0 270.408p 10000.0u 270.409p 0 274.484p 0 274.485p 10000.0u 274.486p 0 289.859p 0 289.86p 10000.0u 289.861p 0 302.138p 0 302.139p 10000.0u 302.14p 0 310.121p 0 310.122p 10000.0u 310.123p 0 315.44p 0 315.441p 10000.0u 315.442p 0 321.92p 0 321.921p 10000.0u 321.922p 0 329.534p 0 329.535p 10000.0u 329.536p 0 335.318p 0 335.319p 10000.0u 335.32p 0 354.224p 0 354.225p 10000.0u 354.226p 0 361.088p 0 361.089p 10000.0u 361.09p 0 362.066p 0 362.067p 10000.0u 362.068p 0 365.171p 0 365.172p 10000.0u 365.173p 0 373.634p 0 373.635p 10000.0u 373.636p 0 399.593p 0 399.594p 10000.0u 399.595p 0 410.786p 0 410.787p 10000.0u 410.788p 0 427.241p 0 427.242p 10000.0u 427.243p 0 441.005p 0 441.006p 10000.0u 441.007p 0 455.354p 0 455.355p 10000.0u 455.356p 0 473.051p 0 473.052p 10000.0u 473.053p 0 473.486p 0 473.487p 10000.0u 473.488p 0 494.318p 0 494.319p 10000.0u 494.32p 0 499.304p 0 499.305p 10000.0u 499.306p 0 500.387p 0 500.388p 10000.0u 500.389p 0 518.321p 0 518.322p 10000.0u 518.323p 0 523.892p 0 523.893p 10000.0u 523.894p 0 528.884p 0 528.885p 10000.0u 528.886p 0 529.358p 0 529.359p 10000.0u 529.36p 0 534.896p 0 534.897p 10000.0u 534.898p 0 550.934p 0 550.935p 10000.0u 550.936p 0 574.541p 0 574.542p 10000.0u 574.543p 0 581.54p 0 581.541p 10000.0u 581.542p 0 593.45p 0 593.451p 10000.0u 593.452p 0 620.126p 0 620.127p 10000.0u 620.128p 0 620.279p 0 620.28p 10000.0u 620.281p 0 631.079p 0 631.08p 10000.0u 631.081p 0 637.652p 0 637.653p 10000.0u 637.654p 0 643.595p 0 643.596p 10000.0u 643.597p 0 674.351p 0 674.352p 10000.0u 674.353p 0 685.463p 0 685.464p 10000.0u 685.465p 0 689.975p 0 689.976p 10000.0u 689.977p 0 704.582p 0 704.583p 10000.0u 704.584p 0 713.873p 0 713.874p 10000.0u 713.875p 0 719.465p 0 719.466p 10000.0u 719.467p 0 742.412p 0 742.413p 10000.0u 742.414p 0 771.53p 0 771.531p 10000.0u 771.532p 0 772.13p 0 772.131p 10000.0u 772.132p 0 785.771p 0 785.772p 10000.0u 785.773p 0 793.415p 0 793.416p 10000.0u 793.417p 0 807.263p 0 807.264p 10000.0u 807.265p 0 820.268p 0 820.269p 10000.0u 820.27p 0 831.989p 0 831.99p 10000.0u 831.991p 0 841.688p 0 841.689p 10000.0u 841.69p 0 849.839p 0 849.84p 10000.0u 849.841p 0 851.36p 0 851.361p 10000.0u 851.362p 0 855.287p 0 855.288p 10000.0u 855.289p 0 866.777p 0 866.778p 10000.0u 866.779p 0 877.994p 0 877.995p 10000.0u 877.996p 0 898.775p 0 898.776p 10000.0u 898.777p 0 909.002p 0 909.003p 10000.0u 909.004p 0 917.414p 0 917.415p 10000.0u 917.416p 0 939.824p 0 939.825p 10000.0u 939.826p 0 948.554p 0 948.555p 10000.0u 948.556p 0 967.61p 0 967.611p 10000.0u 967.612p 0 978.374p 0 978.375p 10000.0u 978.376p 0 982.76p 0 982.761p 10000.0u 982.762p 0 983.078p 0 983.079p 10000.0u 983.08p 0 987.68p 0 987.681p 10000.0u 987.682p 0 988.562p 0 988.563p 10000.0u 988.564p 0 988.703p 0 988.704p 10000.0u 988.705p 0 995.471p 0 995.472p 10000.0u 995.473p 0)
IIN52 0 53 pwl(0 0 1.22p 0 1.221p 10000.0u 1.222p 0 8.537p 0 8.538p 10000.0u 8.539p 0 9.803p 0 9.804p 10000.0u 9.805p 0 11.066p 0 11.067p 10000.0u 11.068p 0 23.645p 0 23.646p 10000.0u 23.647p 0 25.976p 0 25.977p 10000.0u 25.978p 0 49.964p 0 49.965p 10000.0u 49.966p 0 69.005p 0 69.006p 10000.0u 69.007p 0 71.054p 0 71.055p 10000.0u 71.056p 0 76.763p 0 76.764p 10000.0u 76.765p 0 77.681p 0 77.682p 10000.0u 77.683p 0 106.175p 0 106.176p 10000.0u 106.177p 0 128.714p 0 128.715p 10000.0u 128.716p 0 146.324p 0 146.325p 10000.0u 146.326p 0 152.48p 0 152.481p 10000.0u 152.482p 0 167.456p 0 167.457p 10000.0u 167.458p 0 173.657p 0 173.658p 10000.0u 173.659p 0 184.046p 0 184.047p 10000.0u 184.048p 0 201.155p 0 201.156p 10000.0u 201.157p 0 224.42p 0 224.421p 10000.0u 224.422p 0 232.697p 0 232.698p 10000.0u 232.699p 0 266.915p 0 266.916p 10000.0u 266.917p 0 274.394p 0 274.395p 10000.0u 274.396p 0 280.616p 0 280.617p 10000.0u 280.618p 0 289.67p 0 289.671p 10000.0u 289.672p 0 295.589p 0 295.59p 10000.0u 295.591p 0 297.575p 0 297.576p 10000.0u 297.577p 0 314.807p 0 314.808p 10000.0u 314.809p 0 329.234p 0 329.235p 10000.0u 329.236p 0 330.308p 0 330.309p 10000.0u 330.31p 0 356.696p 0 356.697p 10000.0u 356.698p 0 366.599p 0 366.6p 10000.0u 366.601p 0 374.48p 0 374.481p 10000.0u 374.482p 0 387.569p 0 387.57p 10000.0u 387.571p 0 389.252p 0 389.253p 10000.0u 389.254p 0 397.673p 0 397.674p 10000.0u 397.675p 0 414.227p 0 414.228p 10000.0u 414.229p 0 419.195p 0 419.196p 10000.0u 419.197p 0 459.44p 0 459.441p 10000.0u 459.442p 0 462.494p 0 462.495p 10000.0u 462.496p 0 463.904p 0 463.905p 10000.0u 463.906p 0 470.408p 0 470.409p 10000.0u 470.41p 0 478.259p 0 478.26p 10000.0u 478.261p 0 482.186p 0 482.187p 10000.0u 482.188p 0 498.509p 0 498.51p 10000.0u 498.511p 0 502.088p 0 502.089p 10000.0u 502.09p 0 502.574p 0 502.575p 10000.0u 502.576p 0 526.364p 0 526.365p 10000.0u 526.366p 0 532.982p 0 532.983p 10000.0u 532.984p 0 536.546p 0 536.547p 10000.0u 536.548p 0 540.806p 0 540.807p 10000.0u 540.808p 0 557.759p 0 557.76p 10000.0u 557.761p 0 563.309p 0 563.31p 10000.0u 563.311p 0 563.795p 0 563.796p 10000.0u 563.797p 0 579.02p 0 579.021p 10000.0u 579.022p 0 583.901p 0 583.902p 10000.0u 583.903p 0 606.698p 0 606.699p 10000.0u 606.7p 0 611.063p 0 611.064p 10000.0u 611.065p 0 618.194p 0 618.195p 10000.0u 618.196p 0 620.096p 0 620.097p 10000.0u 620.098p 0 634.583p 0 634.584p 10000.0u 634.585p 0 636.512p 0 636.513p 10000.0u 636.514p 0 659.462p 0 659.463p 10000.0u 659.464p 0 669.215p 0 669.216p 10000.0u 669.217p 0 679.106p 0 679.107p 10000.0u 679.108p 0 679.481p 0 679.482p 10000.0u 679.483p 0 692.804p 0 692.805p 10000.0u 692.806p 0 709.193p 0 709.194p 10000.0u 709.195p 0 710.903p 0 710.904p 10000.0u 710.905p 0 712.01p 0 712.011p 10000.0u 712.012p 0 713.624p 0 713.625p 10000.0u 713.626p 0 717.629p 0 717.63p 10000.0u 717.631p 0 721.193p 0 721.194p 10000.0u 721.195p 0 751.604p 0 751.605p 10000.0u 751.606p 0 755.372p 0 755.373p 10000.0u 755.374p 0 756.779p 0 756.78p 10000.0u 756.781p 0 762.527p 0 762.528p 10000.0u 762.529p 0 769.73p 0 769.731p 10000.0u 769.732p 0 777.05p 0 777.051p 10000.0u 777.052p 0 787.472p 0 787.473p 10000.0u 787.474p 0 800.405p 0 800.406p 10000.0u 800.407p 0 817.976p 0 817.977p 10000.0u 817.978p 0 828.893p 0 828.894p 10000.0u 828.895p 0 830.543p 0 830.544p 10000.0u 830.545p 0 835.916p 0 835.917p 10000.0u 835.918p 0 836.651p 0 836.652p 10000.0u 836.653p 0 839.114p 0 839.115p 10000.0u 839.116p 0 854.672p 0 854.673p 10000.0u 854.674p 0 874.349p 0 874.35p 10000.0u 874.351p 0 874.676p 0 874.677p 10000.0u 874.678p 0 882.995p 0 882.996p 10000.0u 882.997p 0 902.975p 0 902.976p 10000.0u 902.977p 0 921.776p 0 921.777p 10000.0u 921.778p 0 929.165p 0 929.166p 10000.0u 929.167p 0 942.497p 0 942.498p 10000.0u 942.499p 0 945.332p 0 945.333p 10000.0u 945.334p 0 945.77p 0 945.771p 10000.0u 945.772p 0 949.97p 0 949.971p 10000.0u 949.972p 0 952.373p 0 952.374p 10000.0u 952.375p 0 964.919p 0 964.92p 10000.0u 964.921p 0 972.293p 0 972.294p 10000.0u 972.295p 0 996.953p 0 996.954p 10000.0u 996.955p 0 997.961p 0 997.962p 10000.0u 997.963p 0)
IIN53 0 54 pwl(0 0 5.078p 0 5.079p 10000.0u 5.08p 0 6.665p 0 6.666p 10000.0u 6.667p 0 8.192p 0 8.193p 10000.0u 8.194p 0 10.049p 0 10.05p 10000.0u 10.051p 0 38.513p 0 38.514p 10000.0u 38.515p 0 44.513p 0 44.514p 10000.0u 44.515p 0 58.85p 0 58.851p 10000.0u 58.852p 0 68.618p 0 68.619p 10000.0u 68.62p 0 99.089p 0 99.09p 10000.0u 99.091p 0 102.947p 0 102.948p 10000.0u 102.949p 0 110.12p 0 110.121p 10000.0u 110.122p 0 113.288p 0 113.289p 10000.0u 113.29p 0 120.884p 0 120.885p 10000.0u 120.886p 0 121.97p 0 121.971p 10000.0u 121.972p 0 137.294p 0 137.295p 10000.0u 137.296p 0 167.642p 0 167.643p 10000.0u 167.644p 0 168.74p 0 168.741p 10000.0u 168.742p 0 183.065p 0 183.066p 10000.0u 183.067p 0 183.272p 0 183.273p 10000.0u 183.274p 0 190.907p 0 190.908p 10000.0u 190.909p 0 195.929p 0 195.93p 10000.0u 195.931p 0 197.042p 0 197.043p 10000.0u 197.044p 0 200.732p 0 200.733p 10000.0u 200.734p 0 205.109p 0 205.11p 10000.0u 205.111p 0 205.778p 0 205.779p 10000.0u 205.78p 0 209.873p 0 209.874p 10000.0u 209.875p 0 225.965p 0 225.966p 10000.0u 225.967p 0 250.922p 0 250.923p 10000.0u 250.924p 0 271.769p 0 271.77p 10000.0u 271.771p 0 276.5p 0 276.501p 10000.0u 276.502p 0 289.706p 0 289.707p 10000.0u 289.708p 0 306.17p 0 306.171p 10000.0u 306.172p 0 310.457p 0 310.458p 10000.0u 310.459p 0 326.846p 0 326.847p 10000.0u 326.848p 0 341.735p 0 341.736p 10000.0u 341.737p 0 356.03p 0 356.031p 10000.0u 356.032p 0 357.125p 0 357.126p 10000.0u 357.127p 0 370.568p 0 370.569p 10000.0u 370.57p 0 372.113p 0 372.114p 10000.0u 372.115p 0 376.451p 0 376.452p 10000.0u 376.453p 0 377.483p 0 377.484p 10000.0u 377.485p 0 378.134p 0 378.135p 10000.0u 378.136p 0 403.67p 0 403.671p 10000.0u 403.672p 0 408.914p 0 408.915p 10000.0u 408.916p 0 413.921p 0 413.922p 10000.0u 413.923p 0 420.524p 0 420.525p 10000.0u 420.526p 0 431.744p 0 431.745p 10000.0u 431.746p 0 478.757p 0 478.758p 10000.0u 478.759p 0 479.006p 0 479.007p 10000.0u 479.008p 0 489.098p 0 489.099p 10000.0u 489.1p 0 499.844p 0 499.845p 10000.0u 499.846p 0 532.952p 0 532.953p 10000.0u 532.954p 0 538.514p 0 538.515p 10000.0u 538.516p 0 541.262p 0 541.263p 10000.0u 541.264p 0 542.606p 0 542.607p 10000.0u 542.608p 0 548.54p 0 548.541p 10000.0u 548.542p 0 576.041p 0 576.042p 10000.0u 576.043p 0 586.808p 0 586.809p 10000.0u 586.81p 0 608.855p 0 608.856p 10000.0u 608.857p 0 609.665p 0 609.666p 10000.0u 609.667p 0 613.196p 0 613.197p 10000.0u 613.198p 0 648.533p 0 648.534p 10000.0u 648.535p 0 650.177p 0 650.178p 10000.0u 650.179p 0 653.987p 0 653.988p 10000.0u 653.989p 0 657.653p 0 657.654p 10000.0u 657.655p 0 684.209p 0 684.21p 10000.0u 684.211p 0 684.365p 0 684.366p 10000.0u 684.367p 0 701.006p 0 701.007p 10000.0u 701.008p 0 708.311p 0 708.312p 10000.0u 708.313p 0 710.516p 0 710.517p 10000.0u 710.518p 0 721.196p 0 721.197p 10000.0u 721.198p 0 723.887p 0 723.888p 10000.0u 723.889p 0 734.507p 0 734.508p 10000.0u 734.509p 0 745.022p 0 745.023p 10000.0u 745.024p 0 751.877p 0 751.878p 10000.0u 751.879p 0 760.727p 0 760.728p 10000.0u 760.729p 0 762.899p 0 762.9p 10000.0u 762.901p 0 766.652p 0 766.653p 10000.0u 766.654p 0 768.812p 0 768.813p 10000.0u 768.814p 0 779.3p 0 779.301p 10000.0u 779.302p 0 794.588p 0 794.589p 10000.0u 794.59p 0 795.587p 0 795.588p 10000.0u 795.589p 0 798.599p 0 798.6p 10000.0u 798.601p 0 804.635p 0 804.636p 10000.0u 804.637p 0 813.161p 0 813.162p 10000.0u 813.163p 0 819.782p 0 819.783p 10000.0u 819.784p 0 871.322p 0 871.323p 10000.0u 871.324p 0 872.807p 0 872.808p 10000.0u 872.809p 0 875.366p 0 875.367p 10000.0u 875.368p 0 877.496p 0 877.497p 10000.0u 877.498p 0 902.225p 0 902.226p 10000.0u 902.227p 0 923.39p 0 923.391p 10000.0u 923.392p 0 930.215p 0 930.216p 10000.0u 930.217p 0 941.573p 0 941.574p 10000.0u 941.575p 0 945.773p 0 945.774p 10000.0u 945.775p 0 950.285p 0 950.286p 10000.0u 950.287p 0 953.477p 0 953.478p 10000.0u 953.479p 0 962.693p 0 962.694p 10000.0u 962.695p 0 968.054p 0 968.055p 10000.0u 968.056p 0 970.988p 0 970.989p 10000.0u 970.99p 0 972.515p 0 972.516p 10000.0u 972.517p 0 975.383p 0 975.384p 10000.0u 975.385p 0 982.583p 0 982.584p 10000.0u 982.585p 0 982.946p 0 982.947p 10000.0u 982.948p 0 988.823p 0 988.824p 10000.0u 988.825p 0 992.957p 0 992.958p 10000.0u 992.959p 0 994.199p 0 994.2p 10000.0u 994.201p 0)
IIN54 0 55 pwl(0 0 14.369p 0 14.37p 10000.0u 14.371p 0 33.218p 0 33.219p 10000.0u 33.22p 0 48.494p 0 48.495p 10000.0u 48.496p 0 56.84p 0 56.841p 10000.0u 56.842p 0 58.946p 0 58.947p 10000.0u 58.948p 0 59.756p 0 59.757p 10000.0u 59.758p 0 62.447p 0 62.448p 10000.0u 62.449p 0 68.711p 0 68.712p 10000.0u 68.713p 0 76.097p 0 76.098p 10000.0u 76.099p 0 99.026p 0 99.027p 10000.0u 99.028p 0 116.114p 0 116.115p 10000.0u 116.116p 0 116.285p 0 116.286p 10000.0u 116.287p 0 116.507p 0 116.508p 10000.0u 116.509p 0 118.637p 0 118.638p 10000.0u 118.639p 0 122.429p 0 122.43p 10000.0u 122.431p 0 139.061p 0 139.062p 10000.0u 139.063p 0 149.042p 0 149.043p 10000.0u 149.044p 0 154.406p 0 154.407p 10000.0u 154.408p 0 158.447p 0 158.448p 10000.0u 158.449p 0 160.028p 0 160.029p 10000.0u 160.03p 0 165.227p 0 165.228p 10000.0u 165.229p 0 165.926p 0 165.927p 10000.0u 165.928p 0 173.771p 0 173.772p 10000.0u 173.773p 0 173.897p 0 173.898p 10000.0u 173.899p 0 181.067p 0 181.068p 10000.0u 181.069p 0 182.294p 0 182.295p 10000.0u 182.296p 0 182.594p 0 182.595p 10000.0u 182.596p 0 203.081p 0 203.082p 10000.0u 203.083p 0 205.808p 0 205.809p 10000.0u 205.81p 0 224.432p 0 224.433p 10000.0u 224.434p 0 265.715p 0 265.716p 10000.0u 265.717p 0 297.833p 0 297.834p 10000.0u 297.835p 0 309.032p 0 309.033p 10000.0u 309.034p 0 310.661p 0 310.662p 10000.0u 310.663p 0 340.118p 0 340.119p 10000.0u 340.12p 0 351.338p 0 351.339p 10000.0u 351.34p 0 351.944p 0 351.945p 10000.0u 351.946p 0 380.696p 0 380.697p 10000.0u 380.698p 0 420.923p 0 420.924p 10000.0u 420.925p 0 423.695p 0 423.696p 10000.0u 423.697p 0 423.938p 0 423.939p 10000.0u 423.94p 0 429.152p 0 429.153p 10000.0u 429.154p 0 435.68p 0 435.681p 10000.0u 435.682p 0 476.483p 0 476.484p 10000.0u 476.485p 0 483.869p 0 483.87p 10000.0u 483.871p 0 487.598p 0 487.599p 10000.0u 487.6p 0 495.797p 0 495.798p 10000.0u 495.799p 0 495.98p 0 495.981p 10000.0u 495.982p 0 510.479p 0 510.48p 10000.0u 510.481p 0 520.301p 0 520.302p 10000.0u 520.303p 0 560.579p 0 560.58p 10000.0u 560.581p 0 576.815p 0 576.816p 10000.0u 576.817p 0 589.901p 0 589.902p 10000.0u 589.903p 0 589.979p 0 589.98p 10000.0u 589.981p 0 590.351p 0 590.352p 10000.0u 590.353p 0 595.316p 0 595.317p 10000.0u 595.318p 0 616.454p 0 616.455p 10000.0u 616.456p 0 631.058p 0 631.059p 10000.0u 631.06p 0 644.948p 0 644.949p 10000.0u 644.95p 0 665.999p 0 666.0p 10000.0u 666.001p 0 686.648p 0 686.649p 10000.0u 686.65p 0 692.855p 0 692.856p 10000.0u 692.857p 0 693.515p 0 693.516p 10000.0u 693.517p 0 698.438p 0 698.439p 10000.0u 698.44p 0 712.322p 0 712.323p 10000.0u 712.324p 0 728.681p 0 728.682p 10000.0u 728.683p 0 761.912p 0 761.913p 10000.0u 761.914p 0 764.018p 0 764.019p 10000.0u 764.02p 0 771.2p 0 771.201p 10000.0u 771.202p 0 771.215p 0 771.216p 10000.0u 771.217p 0 776.444p 0 776.445p 10000.0u 776.446p 0 784.982p 0 784.983p 10000.0u 784.984p 0 788.594p 0 788.595p 10000.0u 788.596p 0 795.683p 0 795.684p 10000.0u 795.685p 0 802.109p 0 802.11p 10000.0u 802.111p 0 815.819p 0 815.82p 10000.0u 815.821p 0 841.325p 0 841.326p 10000.0u 841.327p 0 844.025p 0 844.026p 10000.0u 844.027p 0 857.309p 0 857.31p 10000.0u 857.311p 0 868.166p 0 868.167p 10000.0u 868.168p 0 879.008p 0 879.009p 10000.0u 879.01p 0 912.806p 0 912.807p 10000.0u 912.808p 0 915.254p 0 915.255p 10000.0u 915.256p 0 922.433p 0 922.434p 10000.0u 922.435p 0 959.684p 0 959.685p 10000.0u 959.686p 0 968.63p 0 968.631p 10000.0u 968.632p 0 992.384p 0 992.385p 10000.0u 992.386p 0 994.898p 0 994.899p 10000.0u 994.9p 0)
IIN55 0 56 pwl(0 0 2.708p 0 2.709p 10000.0u 2.71p 0 7.274p 0 7.275p 10000.0u 7.276p 0 12.065p 0 12.066p 10000.0u 12.067p 0 19.766p 0 19.767p 10000.0u 19.768p 0 35.915p 0 35.916p 10000.0u 35.917p 0 40.382p 0 40.383p 10000.0u 40.384p 0 49.28p 0 49.281p 10000.0u 49.282p 0 52.967p 0 52.968p 10000.0u 52.969p 0 65.294p 0 65.295p 10000.0u 65.296p 0 68.264p 0 68.265p 10000.0u 68.266p 0 77.453p 0 77.454p 10000.0u 77.455p 0 88.667p 0 88.668p 10000.0u 88.669p 0 90.743p 0 90.744p 10000.0u 90.745p 0 99.008p 0 99.009p 10000.0u 99.01p 0 106.145p 0 106.146p 10000.0u 106.147p 0 122.387p 0 122.388p 10000.0u 122.389p 0 130.133p 0 130.134p 10000.0u 130.135p 0 133.877p 0 133.878p 10000.0u 133.879p 0 138.533p 0 138.534p 10000.0u 138.535p 0 155.465p 0 155.466p 10000.0u 155.467p 0 166.805p 0 166.806p 10000.0u 166.807p 0 194.972p 0 194.973p 10000.0u 194.974p 0 210.797p 0 210.798p 10000.0u 210.799p 0 213.392p 0 213.393p 10000.0u 213.394p 0 230.549p 0 230.55p 10000.0u 230.551p 0 239.693p 0 239.694p 10000.0u 239.695p 0 248.24p 0 248.241p 10000.0u 248.242p 0 259.601p 0 259.602p 10000.0u 259.603p 0 270.029p 0 270.03p 10000.0u 270.031p 0 284.432p 0 284.433p 10000.0u 284.434p 0 292.682p 0 292.683p 10000.0u 292.684p 0 299.96p 0 299.961p 10000.0u 299.962p 0 306.833p 0 306.834p 10000.0u 306.835p 0 317.414p 0 317.415p 10000.0u 317.416p 0 317.96p 0 317.961p 10000.0u 317.962p 0 332.264p 0 332.265p 10000.0u 332.266p 0 340.694p 0 340.695p 10000.0u 340.696p 0 341.27p 0 341.271p 10000.0u 341.272p 0 348.845p 0 348.846p 10000.0u 348.847p 0 373.778p 0 373.779p 10000.0u 373.78p 0 375.752p 0 375.753p 10000.0u 375.754p 0 380.174p 0 380.175p 10000.0u 380.176p 0 384.515p 0 384.516p 10000.0u 384.517p 0 386.564p 0 386.565p 10000.0u 386.566p 0 406.043p 0 406.044p 10000.0u 406.045p 0 419.696p 0 419.697p 10000.0u 419.698p 0 448.298p 0 448.299p 10000.0u 448.3p 0 456.746p 0 456.747p 10000.0u 456.748p 0 492.002p 0 492.003p 10000.0u 492.004p 0 498.974p 0 498.975p 10000.0u 498.976p 0 505.868p 0 505.869p 10000.0u 505.87p 0 525.635p 0 525.636p 10000.0u 525.637p 0 532.532p 0 532.533p 10000.0u 532.534p 0 550.928p 0 550.929p 10000.0u 550.93p 0 561.773p 0 561.774p 10000.0u 561.775p 0 562.283p 0 562.284p 10000.0u 562.285p 0 569.24p 0 569.241p 10000.0u 569.242p 0 603.143p 0 603.144p 10000.0u 603.145p 0 608.708p 0 608.709p 10000.0u 608.71p 0 620.033p 0 620.034p 10000.0u 620.035p 0 627.929p 0 627.93p 10000.0u 627.931p 0 628.052p 0 628.053p 10000.0u 628.054p 0 645.134p 0 645.135p 10000.0u 645.136p 0 647.846p 0 647.847p 10000.0u 647.848p 0 648.578p 0 648.579p 10000.0u 648.58p 0 648.641p 0 648.642p 10000.0u 648.643p 0 654.518p 0 654.519p 10000.0u 654.52p 0 661.013p 0 661.014p 10000.0u 661.015p 0 664.469p 0 664.47p 10000.0u 664.471p 0 687.482p 0 687.483p 10000.0u 687.484p 0 733.496p 0 733.497p 10000.0u 733.498p 0 761.108p 0 761.109p 10000.0u 761.11p 0 771.896p 0 771.897p 10000.0u 771.898p 0 789.659p 0 789.66p 10000.0u 789.661p 0 789.782p 0 789.783p 10000.0u 789.784p 0 795.482p 0 795.483p 10000.0u 795.484p 0 797.366p 0 797.367p 10000.0u 797.368p 0 802.112p 0 802.113p 10000.0u 802.114p 0 802.67p 0 802.671p 10000.0u 802.672p 0 807.056p 0 807.057p 10000.0u 807.058p 0 812.159p 0 812.16p 10000.0u 812.161p 0 827.678p 0 827.679p 10000.0u 827.68p 0 845.723p 0 845.724p 10000.0u 845.725p 0 872.021p 0 872.022p 10000.0u 872.023p 0 876.47p 0 876.471p 10000.0u 876.472p 0 910.841p 0 910.842p 10000.0u 910.843p 0 936.161p 0 936.162p 10000.0u 936.163p 0 939.131p 0 939.132p 10000.0u 939.133p 0 958.22p 0 958.221p 10000.0u 958.222p 0 958.604p 0 958.605p 10000.0u 958.606p 0 959.018p 0 959.019p 10000.0u 959.02p 0 976.79p 0 976.791p 10000.0u 976.792p 0 979.961p 0 979.962p 10000.0u 979.963p 0)
IIN56 0 57 pwl(0 0 32.501p 0 32.502p 10000.0u 32.503p 0 44.588p 0 44.589p 10000.0u 44.59p 0 66.059p 0 66.06p 10000.0u 66.061p 0 72.794p 0 72.795p 10000.0u 72.796p 0 77.687p 0 77.688p 10000.0u 77.689p 0 79.094p 0 79.095p 10000.0u 79.096p 0 86.282p 0 86.283p 10000.0u 86.284p 0 97.37p 0 97.371p 10000.0u 97.372p 0 102.752p 0 102.753p 10000.0u 102.754p 0 119.567p 0 119.568p 10000.0u 119.569p 0 167.474p 0 167.475p 10000.0u 167.476p 0 173.87p 0 173.871p 10000.0u 173.872p 0 180.386p 0 180.387p 10000.0u 180.388p 0 218.984p 0 218.985p 10000.0u 218.986p 0 219.212p 0 219.213p 10000.0u 219.214p 0 221.978p 0 221.979p 10000.0u 221.98p 0 250.052p 0 250.053p 10000.0u 250.054p 0 251.582p 0 251.583p 10000.0u 251.584p 0 303.347p 0 303.348p 10000.0u 303.349p 0 317.444p 0 317.445p 10000.0u 317.446p 0 327.272p 0 327.273p 10000.0u 327.274p 0 341.285p 0 341.286p 10000.0u 341.287p 0 341.621p 0 341.622p 10000.0u 341.623p 0 350.909p 0 350.91p 10000.0u 350.911p 0 351.851p 0 351.852p 10000.0u 351.853p 0 355.22p 0 355.221p 10000.0u 355.222p 0 363.17p 0 363.171p 10000.0u 363.172p 0 371.255p 0 371.256p 10000.0u 371.257p 0 380.585p 0 380.586p 10000.0u 380.587p 0 397.376p 0 397.377p 10000.0u 397.378p 0 404.243p 0 404.244p 10000.0u 404.245p 0 407.528p 0 407.529p 10000.0u 407.53p 0 422.066p 0 422.067p 10000.0u 422.068p 0 424.649p 0 424.65p 10000.0u 424.651p 0 454.208p 0 454.209p 10000.0u 454.21p 0 458.027p 0 458.028p 10000.0u 458.029p 0 471.863p 0 471.864p 10000.0u 471.865p 0 479.678p 0 479.679p 10000.0u 479.68p 0 509.456p 0 509.457p 10000.0u 509.458p 0 510.194p 0 510.195p 10000.0u 510.196p 0 512.879p 0 512.88p 10000.0u 512.881p 0 515.738p 0 515.739p 10000.0u 515.74p 0 547.892p 0 547.893p 10000.0u 547.894p 0 563.879p 0 563.88p 10000.0u 563.881p 0 564.182p 0 564.183p 10000.0u 564.184p 0 565.643p 0 565.644p 10000.0u 565.645p 0 567.536p 0 567.537p 10000.0u 567.538p 0 580.232p 0 580.233p 10000.0u 580.234p 0 581.897p 0 581.898p 10000.0u 581.899p 0 590.69p 0 590.691p 10000.0u 590.692p 0 595.526p 0 595.527p 10000.0u 595.528p 0 627.05p 0 627.051p 10000.0u 627.052p 0 653.999p 0 654.0p 10000.0u 654.001p 0 680.684p 0 680.685p 10000.0u 680.686p 0 708.674p 0 708.675p 10000.0u 708.676p 0 714.161p 0 714.162p 10000.0u 714.163p 0 720.752p 0 720.753p 10000.0u 720.754p 0 725.231p 0 725.232p 10000.0u 725.233p 0 726.998p 0 726.999p 10000.0u 727.0p 0 736.286p 0 736.287p 10000.0u 736.288p 0 742.946p 0 742.947p 10000.0u 742.948p 0 745.106p 0 745.107p 10000.0u 745.108p 0 747.422p 0 747.423p 10000.0u 747.424p 0 759.788p 0 759.789p 10000.0u 759.79p 0 765.44p 0 765.441p 10000.0u 765.442p 0 765.449p 0 765.45p 10000.0u 765.451p 0 773.495p 0 773.496p 10000.0u 773.497p 0 778.469p 0 778.47p 10000.0u 778.471p 0 785.291p 0 785.292p 10000.0u 785.293p 0 794.723p 0 794.724p 10000.0u 794.725p 0 797.885p 0 797.886p 10000.0u 797.887p 0 811.973p 0 811.974p 10000.0u 811.975p 0 813.071p 0 813.072p 10000.0u 813.073p 0 816.632p 0 816.633p 10000.0u 816.634p 0 826.283p 0 826.284p 10000.0u 826.285p 0 830.801p 0 830.802p 10000.0u 830.803p 0 841.982p 0 841.983p 10000.0u 841.984p 0 846.245p 0 846.246p 10000.0u 846.247p 0 847.175p 0 847.176p 10000.0u 847.177p 0 857.126p 0 857.127p 10000.0u 857.128p 0 862.457p 0 862.458p 10000.0u 862.459p 0 874.886p 0 874.887p 10000.0u 874.888p 0 894.224p 0 894.225p 10000.0u 894.226p 0 899.663p 0 899.664p 10000.0u 899.665p 0 901.355p 0 901.356p 10000.0u 901.357p 0 919.421p 0 919.422p 10000.0u 919.423p 0 952.34p 0 952.341p 10000.0u 952.342p 0 952.706p 0 952.707p 10000.0u 952.708p 0 958.79p 0 958.791p 10000.0u 958.792p 0 963.893p 0 963.894p 10000.0u 963.895p 0 964.049p 0 964.05p 10000.0u 964.051p 0 964.808p 0 964.809p 10000.0u 964.81p 0 970.238p 0 970.239p 10000.0u 970.24p 0 988.733p 0 988.734p 10000.0u 988.735p 0)
IIN57 0 58 pwl(0 0 18.497p 0 18.498p 10000.0u 18.499p 0 22.373p 0 22.374p 10000.0u 22.375p 0 30.41p 0 30.411p 10000.0u 30.412p 0 40.964p 0 40.965p 10000.0u 40.966p 0 55.814p 0 55.815p 10000.0u 55.816p 0 66.146p 0 66.147p 10000.0u 66.148p 0 79.937p 0 79.938p 10000.0u 79.939p 0 103.613p 0 103.614p 10000.0u 103.615p 0 133.919p 0 133.92p 10000.0u 133.921p 0 181.43p 0 181.431p 10000.0u 181.432p 0 187.172p 0 187.173p 10000.0u 187.174p 0 221.228p 0 221.229p 10000.0u 221.23p 0 223.634p 0 223.635p 10000.0u 223.636p 0 240.881p 0 240.882p 10000.0u 240.883p 0 241.253p 0 241.254p 10000.0u 241.255p 0 248.93p 0 248.931p 10000.0u 248.932p 0 254.606p 0 254.607p 10000.0u 254.608p 0 286.022p 0 286.023p 10000.0u 286.024p 0 339.851p 0 339.852p 10000.0u 339.853p 0 346.481p 0 346.482p 10000.0u 346.483p 0 348.908p 0 348.909p 10000.0u 348.91p 0 352.559p 0 352.56p 10000.0u 352.561p 0 369.191p 0 369.192p 10000.0u 369.193p 0 400.532p 0 400.533p 10000.0u 400.534p 0 401.789p 0 401.79p 10000.0u 401.791p 0 429.272p 0 429.273p 10000.0u 429.274p 0 441.794p 0 441.795p 10000.0u 441.796p 0 500.891p 0 500.892p 10000.0u 500.893p 0 503.09p 0 503.091p 10000.0u 503.092p 0 505.478p 0 505.479p 10000.0u 505.48p 0 506.174p 0 506.175p 10000.0u 506.176p 0 512.462p 0 512.463p 10000.0u 512.464p 0 528.689p 0 528.69p 10000.0u 528.691p 0 538.703p 0 538.704p 10000.0u 538.705p 0 555.494p 0 555.495p 10000.0u 555.496p 0 556.559p 0 556.56p 10000.0u 556.561p 0 576.431p 0 576.432p 10000.0u 576.433p 0 594.236p 0 594.237p 10000.0u 594.238p 0 595.532p 0 595.533p 10000.0u 595.534p 0 628.364p 0 628.365p 10000.0u 628.366p 0 630.059p 0 630.06p 10000.0u 630.061p 0 641.063p 0 641.064p 10000.0u 641.065p 0 642.242p 0 642.243p 10000.0u 642.244p 0 646.595p 0 646.596p 10000.0u 646.597p 0 665.474p 0 665.475p 10000.0u 665.476p 0 665.594p 0 665.595p 10000.0u 665.596p 0 672.452p 0 672.453p 10000.0u 672.454p 0 695.624p 0 695.625p 10000.0u 695.626p 0 699.416p 0 699.417p 10000.0u 699.418p 0 703.013p 0 703.014p 10000.0u 703.015p 0 708.263p 0 708.264p 10000.0u 708.265p 0 711.302p 0 711.303p 10000.0u 711.304p 0 722.435p 0 722.436p 10000.0u 722.437p 0 734.435p 0 734.436p 10000.0u 734.437p 0 735.377p 0 735.378p 10000.0u 735.379p 0 743.093p 0 743.094p 10000.0u 743.095p 0 746.972p 0 746.973p 10000.0u 746.974p 0 769.289p 0 769.29p 10000.0u 769.291p 0 780.599p 0 780.6p 10000.0u 780.601p 0 791.375p 0 791.376p 10000.0u 791.377p 0 795.773p 0 795.774p 10000.0u 795.775p 0 802.004p 0 802.005p 10000.0u 802.006p 0 802.46p 0 802.461p 10000.0u 802.462p 0 814.109p 0 814.11p 10000.0u 814.111p 0 843.293p 0 843.294p 10000.0u 843.295p 0 868.673p 0 868.674p 10000.0u 868.675p 0 877.613p 0 877.614p 10000.0u 877.615p 0 935.072p 0 935.073p 10000.0u 935.074p 0 949.727p 0 949.728p 10000.0u 949.729p 0 990.725p 0 990.726p 10000.0u 990.727p 0 992.498p 0 992.499p 10000.0u 992.5p 0)
IIN58 0 59 pwl(0 0 0.998p 0 0.999p 10000.0u 1.0p 0 25.265p 0 25.266p 10000.0u 25.267p 0 41.531p 0 41.532p 10000.0u 41.533p 0 52.109p 0 52.11p 10000.0u 52.111p 0 70.556p 0 70.557p 10000.0u 70.558p 0 70.631p 0 70.632p 10000.0u 70.633p 0 78.074p 0 78.075p 10000.0u 78.076p 0 86.528p 0 86.529p 10000.0u 86.53p 0 105.743p 0 105.744p 10000.0u 105.745p 0 106.997p 0 106.998p 10000.0u 106.999p 0 129.689p 0 129.69p 10000.0u 129.691p 0 167.639p 0 167.64p 10000.0u 167.641p 0 176.564p 0 176.565p 10000.0u 176.566p 0 177.377p 0 177.378p 10000.0u 177.379p 0 185.792p 0 185.793p 10000.0u 185.794p 0 191.9p 0 191.901p 10000.0u 191.902p 0 214.799p 0 214.8p 10000.0u 214.801p 0 224.015p 0 224.016p 10000.0u 224.017p 0 235.178p 0 235.179p 10000.0u 235.18p 0 241.274p 0 241.275p 10000.0u 241.276p 0 253.466p 0 253.467p 10000.0u 253.468p 0 259.511p 0 259.512p 10000.0u 259.513p 0 285.878p 0 285.879p 10000.0u 285.88p 0 292.859p 0 292.86p 10000.0u 292.861p 0 293.402p 0 293.403p 10000.0u 293.404p 0 296.939p 0 296.94p 10000.0u 296.941p 0 297.803p 0 297.804p 10000.0u 297.805p 0 297.806p 0 297.807p 10000.0u 297.808p 0 300.734p 0 300.735p 10000.0u 300.736p 0 301.583p 0 301.584p 10000.0u 301.585p 0 301.913p 0 301.914p 10000.0u 301.915p 0 302.753p 0 302.754p 10000.0u 302.755p 0 307.127p 0 307.128p 10000.0u 307.129p 0 336.077p 0 336.078p 10000.0u 336.079p 0 341.828p 0 341.829p 10000.0u 341.83p 0 341.918p 0 341.919p 10000.0u 341.92p 0 345.155p 0 345.156p 10000.0u 345.157p 0 373.958p 0 373.959p 10000.0u 373.96p 0 413.84p 0 413.841p 10000.0u 413.842p 0 438.11p 0 438.111p 10000.0u 438.112p 0 483.47p 0 483.471p 10000.0u 483.472p 0 490.199p 0 490.2p 10000.0u 490.201p 0 512.828p 0 512.829p 10000.0u 512.83p 0 527.786p 0 527.787p 10000.0u 527.788p 0 545.219p 0 545.22p 10000.0u 545.221p 0 546.38p 0 546.381p 10000.0u 546.382p 0 549.179p 0 549.18p 10000.0u 549.181p 0 589.766p 0 589.767p 10000.0u 589.768p 0 590.777p 0 590.778p 10000.0u 590.779p 0 597.047p 0 597.048p 10000.0u 597.049p 0 598.856p 0 598.857p 10000.0u 598.858p 0 606.17p 0 606.171p 10000.0u 606.172p 0 616.049p 0 616.05p 10000.0u 616.051p 0 622.637p 0 622.638p 10000.0u 622.639p 0 624.326p 0 624.327p 10000.0u 624.328p 0 625.316p 0 625.317p 10000.0u 625.318p 0 658.373p 0 658.374p 10000.0u 658.375p 0 682.556p 0 682.557p 10000.0u 682.558p 0 685.604p 0 685.605p 10000.0u 685.606p 0 694.907p 0 694.908p 10000.0u 694.909p 0 719.627p 0 719.628p 10000.0u 719.629p 0 755.912p 0 755.913p 10000.0u 755.914p 0 762.221p 0 762.222p 10000.0u 762.223p 0 768.011p 0 768.012p 10000.0u 768.013p 0 777.176p 0 777.177p 10000.0u 777.178p 0 778.067p 0 778.068p 10000.0u 778.069p 0 798.455p 0 798.456p 10000.0u 798.457p 0 806.969p 0 806.97p 10000.0u 806.971p 0 807.608p 0 807.609p 10000.0u 807.61p 0 812.207p 0 812.208p 10000.0u 812.209p 0 815.528p 0 815.529p 10000.0u 815.53p 0 824.525p 0 824.526p 10000.0u 824.527p 0 835.079p 0 835.08p 10000.0u 835.081p 0 860.294p 0 860.295p 10000.0u 860.296p 0 867.152p 0 867.153p 10000.0u 867.154p 0 885.587p 0 885.588p 10000.0u 885.589p 0 891.659p 0 891.66p 10000.0u 891.661p 0 927.362p 0 927.363p 10000.0u 927.364p 0 931.445p 0 931.446p 10000.0u 931.447p 0 951.965p 0 951.966p 10000.0u 951.967p 0 959.915p 0 959.916p 10000.0u 959.917p 0 965.006p 0 965.007p 10000.0u 965.008p 0 973.964p 0 973.965p 10000.0u 973.966p 0 977.486p 0 977.487p 10000.0u 977.488p 0 980.363p 0 980.364p 10000.0u 980.365p 0 985.436p 0 985.437p 10000.0u 985.438p 0 991.277p 0 991.278p 10000.0u 991.279p 0 996.02p 0 996.021p 10000.0u 996.022p 0 998.141p 0 998.142p 10000.0u 998.143p 0)
IIN59 0 60 pwl(0 0 15.587p 0 15.588p 10000.0u 15.589p 0 19.976p 0 19.977p 10000.0u 19.978p 0 24.869p 0 24.87p 10000.0u 24.871p 0 38.174p 0 38.175p 10000.0u 38.176p 0 40.016p 0 40.017p 10000.0u 40.018p 0 50.477p 0 50.478p 10000.0u 50.479p 0 52.994p 0 52.995p 10000.0u 52.996p 0 62.318p 0 62.319p 10000.0u 62.32p 0 63.275p 0 63.276p 10000.0u 63.277p 0 94.481p 0 94.482p 10000.0u 94.483p 0 104.909p 0 104.91p 10000.0u 104.911p 0 106.103p 0 106.104p 10000.0u 106.105p 0 135.374p 0 135.375p 10000.0u 135.376p 0 146.498p 0 146.499p 10000.0u 146.5p 0 155.597p 0 155.598p 10000.0u 155.599p 0 184.487p 0 184.488p 10000.0u 184.489p 0 194.297p 0 194.298p 10000.0u 194.299p 0 194.996p 0 194.997p 10000.0u 194.998p 0 208.769p 0 208.77p 10000.0u 208.771p 0 210.746p 0 210.747p 10000.0u 210.748p 0 216.803p 0 216.804p 10000.0u 216.805p 0 221.699p 0 221.7p 10000.0u 221.701p 0 221.972p 0 221.973p 10000.0u 221.974p 0 239.597p 0 239.598p 10000.0u 239.599p 0 242.066p 0 242.067p 10000.0u 242.068p 0 251.711p 0 251.712p 10000.0u 251.713p 0 251.813p 0 251.814p 10000.0u 251.815p 0 278.369p 0 278.37p 10000.0u 278.371p 0 282.884p 0 282.885p 10000.0u 282.886p 0 290.255p 0 290.256p 10000.0u 290.257p 0 300.428p 0 300.429p 10000.0u 300.43p 0 305.663p 0 305.664p 10000.0u 305.665p 0 313.265p 0 313.266p 10000.0u 313.267p 0 329.405p 0 329.406p 10000.0u 329.407p 0 340.127p 0 340.128p 10000.0u 340.129p 0 343.895p 0 343.896p 10000.0u 343.897p 0 344.75p 0 344.751p 10000.0u 344.752p 0 373.715p 0 373.716p 10000.0u 373.717p 0 376.43p 0 376.431p 10000.0u 376.432p 0 403.631p 0 403.632p 10000.0u 403.633p 0 404.438p 0 404.439p 10000.0u 404.44p 0 406.346p 0 406.347p 10000.0u 406.348p 0 424.466p 0 424.467p 10000.0u 424.468p 0 442.007p 0 442.008p 10000.0u 442.009p 0 443.498p 0 443.499p 10000.0u 443.5p 0 450.746p 0 450.747p 10000.0u 450.748p 0 477.2p 0 477.201p 10000.0u 477.202p 0 493.481p 0 493.482p 10000.0u 493.483p 0 506.3p 0 506.301p 10000.0u 506.302p 0 530.273p 0 530.274p 10000.0u 530.275p 0 579.086p 0 579.087p 10000.0u 579.088p 0 583.334p 0 583.335p 10000.0u 583.336p 0 583.628p 0 583.629p 10000.0u 583.63p 0 586.547p 0 586.548p 10000.0u 586.549p 0 588.494p 0 588.495p 10000.0u 588.496p 0 601.463p 0 601.464p 10000.0u 601.465p 0 613.178p 0 613.179p 10000.0u 613.18p 0 649.448p 0 649.449p 10000.0u 649.45p 0 651.788p 0 651.789p 10000.0u 651.79p 0 652.643p 0 652.644p 10000.0u 652.645p 0 656.003p 0 656.004p 10000.0u 656.005p 0 667.517p 0 667.518p 10000.0u 667.519p 0 701.354p 0 701.355p 10000.0u 701.356p 0 704.318p 0 704.319p 10000.0u 704.32p 0 706.943p 0 706.944p 10000.0u 706.945p 0 710.366p 0 710.367p 10000.0u 710.368p 0 733.346p 0 733.347p 10000.0u 733.348p 0 733.505p 0 733.506p 10000.0u 733.507p 0 767.876p 0 767.877p 10000.0u 767.878p 0 768.023p 0 768.024p 10000.0u 768.025p 0 771.89p 0 771.891p 10000.0u 771.892p 0 774.677p 0 774.678p 10000.0u 774.679p 0 774.698p 0 774.699p 10000.0u 774.7p 0 804.341p 0 804.342p 10000.0u 804.343p 0 811.748p 0 811.749p 10000.0u 811.75p 0 815.633p 0 815.634p 10000.0u 815.635p 0 815.699p 0 815.7p 10000.0u 815.701p 0 819.497p 0 819.498p 10000.0u 819.499p 0 824.54p 0 824.541p 10000.0u 824.542p 0 831.524p 0 831.525p 10000.0u 831.526p 0 849.188p 0 849.189p 10000.0u 849.19p 0 851.87p 0 851.871p 10000.0u 851.872p 0 862.319p 0 862.32p 10000.0u 862.321p 0 867.929p 0 867.93p 10000.0u 867.931p 0 876.482p 0 876.483p 10000.0u 876.484p 0 883.253p 0 883.254p 10000.0u 883.255p 0 883.646p 0 883.647p 10000.0u 883.648p 0 887.987p 0 887.988p 10000.0u 887.989p 0 895.04p 0 895.041p 10000.0u 895.042p 0 909.737p 0 909.738p 10000.0u 909.739p 0 909.971p 0 909.972p 10000.0u 909.973p 0 916.958p 0 916.959p 10000.0u 916.96p 0 920.234p 0 920.235p 10000.0u 920.236p 0 934.316p 0 934.317p 10000.0u 934.318p 0 956.162p 0 956.163p 10000.0u 956.164p 0 965.027p 0 965.028p 10000.0u 965.029p 0 968.999p 0 969.0p 10000.0u 969.001p 0 991.181p 0 991.182p 10000.0u 991.183p 0)
IIN60 0 61 pwl(0 0 1.733p 0 1.734p 10000.0u 1.735p 0 6.53p 0 6.531p 10000.0u 6.532p 0 16.697p 0 16.698p 10000.0u 16.699p 0 18.326p 0 18.327p 10000.0u 18.328p 0 27.605p 0 27.606p 10000.0u 27.607p 0 28.676p 0 28.677p 10000.0u 28.678p 0 55.379p 0 55.38p 10000.0u 55.381p 0 75.509p 0 75.51p 10000.0u 75.511p 0 90.83p 0 90.831p 10000.0u 90.832p 0 97.049p 0 97.05p 10000.0u 97.051p 0 109.427p 0 109.428p 10000.0u 109.429p 0 129.47p 0 129.471p 10000.0u 129.472p 0 139.595p 0 139.596p 10000.0u 139.597p 0 150.404p 0 150.405p 10000.0u 150.406p 0 153.137p 0 153.138p 10000.0u 153.139p 0 158.423p 0 158.424p 10000.0u 158.425p 0 183.332p 0 183.333p 10000.0u 183.334p 0 188.564p 0 188.565p 10000.0u 188.566p 0 198.392p 0 198.393p 10000.0u 198.394p 0 212.504p 0 212.505p 10000.0u 212.506p 0 213.443p 0 213.444p 10000.0u 213.445p 0 220.859p 0 220.86p 10000.0u 220.861p 0 224.951p 0 224.952p 10000.0u 224.953p 0 232.604p 0 232.605p 10000.0u 232.606p 0 276.566p 0 276.567p 10000.0u 276.568p 0 278.0p 0 278.001p 10000.0u 278.002p 0 278.165p 0 278.166p 10000.0u 278.167p 0 291.917p 0 291.918p 10000.0u 291.919p 0 312.224p 0 312.225p 10000.0u 312.226p 0 313.271p 0 313.272p 10000.0u 313.273p 0 319.058p 0 319.059p 10000.0u 319.06p 0 348.125p 0 348.126p 10000.0u 348.127p 0 348.371p 0 348.372p 10000.0u 348.373p 0 357.911p 0 357.912p 10000.0u 357.913p 0 367.661p 0 367.662p 10000.0u 367.663p 0 387.077p 0 387.078p 10000.0u 387.079p 0 394.301p 0 394.302p 10000.0u 394.303p 0 394.517p 0 394.518p 10000.0u 394.519p 0 411.572p 0 411.573p 10000.0u 411.574p 0 418.127p 0 418.128p 10000.0u 418.129p 0 436.415p 0 436.416p 10000.0u 436.417p 0 440.774p 0 440.775p 10000.0u 440.776p 0 445.496p 0 445.497p 10000.0u 445.498p 0 448.496p 0 448.497p 10000.0u 448.498p 0 450.461p 0 450.462p 10000.0u 450.463p 0 465.593p 0 465.594p 10000.0u 465.595p 0 465.755p 0 465.756p 10000.0u 465.757p 0 467.237p 0 467.238p 10000.0u 467.239p 0 480.938p 0 480.939p 10000.0u 480.94p 0 482.012p 0 482.013p 10000.0u 482.014p 0 482.255p 0 482.256p 10000.0u 482.257p 0 502.064p 0 502.065p 10000.0u 502.066p 0 502.685p 0 502.686p 10000.0u 502.687p 0 531.779p 0 531.78p 10000.0u 531.781p 0 533.333p 0 533.334p 10000.0u 533.335p 0 536.9p 0 536.901p 10000.0u 536.902p 0 550.817p 0 550.818p 10000.0u 550.819p 0 557.396p 0 557.397p 10000.0u 557.398p 0 558.113p 0 558.114p 10000.0u 558.115p 0 560.123p 0 560.124p 10000.0u 560.125p 0 562.07p 0 562.071p 10000.0u 562.072p 0 567.872p 0 567.873p 10000.0u 567.874p 0 569.432p 0 569.433p 10000.0u 569.434p 0 572.6p 0 572.601p 10000.0u 572.602p 0 574.694p 0 574.695p 10000.0u 574.696p 0 583.445p 0 583.446p 10000.0u 583.447p 0 583.982p 0 583.983p 10000.0u 583.984p 0 592.877p 0 592.878p 10000.0u 592.879p 0 597.047p 0 597.048p 10000.0u 597.049p 0 607.448p 0 607.449p 10000.0u 607.45p 0 628.01p 0 628.011p 10000.0u 628.012p 0 628.796p 0 628.797p 10000.0u 628.798p 0 637.481p 0 637.482p 10000.0u 637.483p 0 658.805p 0 658.806p 10000.0u 658.807p 0 667.838p 0 667.839p 10000.0u 667.84p 0 669.539p 0 669.54p 10000.0u 669.541p 0 691.775p 0 691.776p 10000.0u 691.777p 0 708.983p 0 708.984p 10000.0u 708.985p 0 710.501p 0 710.502p 10000.0u 710.503p 0 714.338p 0 714.339p 10000.0u 714.34p 0 716.66p 0 716.661p 10000.0u 716.662p 0 722.978p 0 722.979p 10000.0u 722.98p 0 750.218p 0 750.219p 10000.0u 750.22p 0 754.781p 0 754.782p 10000.0u 754.783p 0 779.405p 0 779.406p 10000.0u 779.407p 0 806.747p 0 806.748p 10000.0u 806.749p 0 821.621p 0 821.622p 10000.0u 821.623p 0 834.56p 0 834.561p 10000.0u 834.562p 0 836.204p 0 836.205p 10000.0u 836.206p 0 837.545p 0 837.546p 10000.0u 837.547p 0 846.071p 0 846.072p 10000.0u 846.073p 0 856.316p 0 856.317p 10000.0u 856.318p 0 860.876p 0 860.877p 10000.0u 860.878p 0 907.511p 0 907.512p 10000.0u 907.513p 0 928.256p 0 928.257p 10000.0u 928.258p 0 931.577p 0 931.578p 10000.0u 931.579p 0 939.473p 0 939.474p 10000.0u 939.475p 0 939.902p 0 939.903p 10000.0u 939.904p 0 948.074p 0 948.075p 10000.0u 948.076p 0 949.052p 0 949.053p 10000.0u 949.054p 0 959.912p 0 959.913p 10000.0u 959.914p 0 962.387p 0 962.388p 10000.0u 962.389p 0)
IIN61 0 62 pwl(0 0 11.405p 0 11.406p 10000.0u 11.407p 0 26.606p 0 26.607p 10000.0u 26.608p 0 43.424p 0 43.425p 10000.0u 43.426p 0 76.529p 0 76.53p 10000.0u 76.531p 0 86.483p 0 86.484p 10000.0u 86.485p 0 88.412p 0 88.413p 10000.0u 88.414p 0 112.184p 0 112.185p 10000.0u 112.186p 0 118.883p 0 118.884p 10000.0u 118.885p 0 124.313p 0 124.314p 10000.0u 124.315p 0 128.438p 0 128.439p 10000.0u 128.44p 0 133.892p 0 133.893p 10000.0u 133.894p 0 136.19p 0 136.191p 10000.0u 136.192p 0 151.454p 0 151.455p 10000.0u 151.456p 0 155.969p 0 155.97p 10000.0u 155.971p 0 157.547p 0 157.548p 10000.0u 157.549p 0 157.886p 0 157.887p 10000.0u 157.888p 0 169.952p 0 169.953p 10000.0u 169.954p 0 173.225p 0 173.226p 10000.0u 173.227p 0 224.906p 0 224.907p 10000.0u 224.908p 0 228.698p 0 228.699p 10000.0u 228.7p 0 250.985p 0 250.986p 10000.0u 250.987p 0 252.575p 0 252.576p 10000.0u 252.577p 0 254.732p 0 254.733p 10000.0u 254.734p 0 256.097p 0 256.098p 10000.0u 256.099p 0 265.406p 0 265.407p 10000.0u 265.408p 0 268.487p 0 268.488p 10000.0u 268.489p 0 307.217p 0 307.218p 10000.0u 307.219p 0 325.079p 0 325.08p 10000.0u 325.081p 0 335.003p 0 335.004p 10000.0u 335.005p 0 344.822p 0 344.823p 10000.0u 344.824p 0 347.126p 0 347.127p 10000.0u 347.128p 0 352.061p 0 352.062p 10000.0u 352.063p 0 362.402p 0 362.403p 10000.0u 362.404p 0 369.269p 0 369.27p 10000.0u 369.271p 0 372.086p 0 372.087p 10000.0u 372.088p 0 381.731p 0 381.732p 10000.0u 381.733p 0 382.004p 0 382.005p 10000.0u 382.006p 0 384.695p 0 384.696p 10000.0u 384.697p 0 396.422p 0 396.423p 10000.0u 396.424p 0 399.23p 0 399.231p 10000.0u 399.232p 0 407.411p 0 407.412p 10000.0u 407.413p 0 411.707p 0 411.708p 10000.0u 411.709p 0 427.448p 0 427.449p 10000.0u 427.45p 0 437.642p 0 437.643p 10000.0u 437.644p 0 438.425p 0 438.426p 10000.0u 438.427p 0 459.488p 0 459.489p 10000.0u 459.49p 0 477.974p 0 477.975p 10000.0u 477.976p 0 503.735p 0 503.736p 10000.0u 503.737p 0 511.4p 0 511.401p 10000.0u 511.402p 0 512.216p 0 512.217p 10000.0u 512.218p 0 512.837p 0 512.838p 10000.0u 512.839p 0 513.095p 0 513.096p 10000.0u 513.097p 0 529.199p 0 529.2p 10000.0u 529.201p 0 536.567p 0 536.568p 10000.0u 536.569p 0 538.196p 0 538.197p 10000.0u 538.198p 0 544.976p 0 544.977p 10000.0u 544.978p 0 549.905p 0 549.906p 10000.0u 549.907p 0 558.029p 0 558.03p 10000.0u 558.031p 0 558.038p 0 558.039p 10000.0u 558.04p 0 562.352p 0 562.353p 10000.0u 562.354p 0 575.024p 0 575.025p 10000.0u 575.026p 0 578.573p 0 578.574p 10000.0u 578.575p 0 582.761p 0 582.762p 10000.0u 582.763p 0 584.465p 0 584.466p 10000.0u 584.467p 0 591.119p 0 591.12p 10000.0u 591.121p 0 614.3p 0 614.301p 10000.0u 614.302p 0 630.815p 0 630.816p 10000.0u 630.817p 0 663.821p 0 663.822p 10000.0u 663.823p 0 671.966p 0 671.967p 10000.0u 671.968p 0 676.283p 0 676.284p 10000.0u 676.285p 0 685.118p 0 685.119p 10000.0u 685.12p 0 695.558p 0 695.559p 10000.0u 695.56p 0 732.89p 0 732.891p 10000.0u 732.892p 0 741.824p 0 741.825p 10000.0u 741.826p 0 745.445p 0 745.446p 10000.0u 745.447p 0 749.141p 0 749.142p 10000.0u 749.143p 0 755.453p 0 755.454p 10000.0u 755.455p 0 757.205p 0 757.206p 10000.0u 757.207p 0 758.651p 0 758.652p 10000.0u 758.653p 0 759.134p 0 759.135p 10000.0u 759.136p 0 772.328p 0 772.329p 10000.0u 772.33p 0 784.439p 0 784.44p 10000.0u 784.441p 0 793.112p 0 793.113p 10000.0u 793.114p 0 793.751p 0 793.752p 10000.0u 793.753p 0 796.265p 0 796.266p 10000.0u 796.267p 0 797.09p 0 797.091p 10000.0u 797.092p 0 807.857p 0 807.858p 10000.0u 807.859p 0 824.798p 0 824.799p 10000.0u 824.8p 0 831.971p 0 831.972p 10000.0u 831.973p 0 832.67p 0 832.671p 10000.0u 832.672p 0 841.523p 0 841.524p 10000.0u 841.525p 0 846.452p 0 846.453p 10000.0u 846.454p 0 853.52p 0 853.521p 10000.0u 853.522p 0 861.158p 0 861.159p 10000.0u 861.16p 0 866.705p 0 866.706p 10000.0u 866.707p 0 869.249p 0 869.25p 10000.0u 869.251p 0 882.812p 0 882.813p 10000.0u 882.814p 0 892.256p 0 892.257p 10000.0u 892.258p 0 902.462p 0 902.463p 10000.0u 902.464p 0 919.481p 0 919.482p 10000.0u 919.483p 0 958.775p 0 958.776p 10000.0u 958.777p 0 961.787p 0 961.788p 10000.0u 961.789p 0 967.388p 0 967.389p 10000.0u 967.39p 0 984.542p 0 984.543p 10000.0u 984.544p 0 989.456p 0 989.457p 10000.0u 989.458p 0)
IIN62 0 63 pwl(0 0 5.045p 0 5.046p 10000.0u 5.047p 0 14.981p 0 14.982p 10000.0u 14.983p 0 16.202p 0 16.203p 10000.0u 16.204p 0 32.099p 0 32.1p 10000.0u 32.101p 0 38.519p 0 38.52p 10000.0u 38.521p 0 39.542p 0 39.543p 10000.0u 39.544p 0 44.516p 0 44.517p 10000.0u 44.518p 0 48.131p 0 48.132p 10000.0u 48.133p 0 60.206p 0 60.207p 10000.0u 60.208p 0 74.3p 0 74.301p 10000.0u 74.302p 0 75.662p 0 75.663p 10000.0u 75.664p 0 76.604p 0 76.605p 10000.0u 76.606p 0 82.073p 0 82.074p 10000.0u 82.075p 0 103.973p 0 103.974p 10000.0u 103.975p 0 105.293p 0 105.294p 10000.0u 105.295p 0 109.262p 0 109.263p 10000.0u 109.264p 0 113.003p 0 113.004p 10000.0u 113.005p 0 116.546p 0 116.547p 10000.0u 116.548p 0 119.87p 0 119.871p 10000.0u 119.872p 0 137.834p 0 137.835p 10000.0u 137.836p 0 143.072p 0 143.073p 10000.0u 143.074p 0 143.207p 0 143.208p 10000.0u 143.209p 0 149.387p 0 149.388p 10000.0u 149.389p 0 159.854p 0 159.855p 10000.0u 159.856p 0 168.014p 0 168.015p 10000.0u 168.016p 0 201.578p 0 201.579p 10000.0u 201.58p 0 202.904p 0 202.905p 10000.0u 202.906p 0 221.972p 0 221.973p 10000.0u 221.974p 0 227.465p 0 227.466p 10000.0u 227.467p 0 253.166p 0 253.167p 10000.0u 253.168p 0 265.331p 0 265.332p 10000.0u 265.333p 0 265.976p 0 265.977p 10000.0u 265.978p 0 269.471p 0 269.472p 10000.0u 269.473p 0 276.194p 0 276.195p 10000.0u 276.196p 0 284.504p 0 284.505p 10000.0u 284.506p 0 300.914p 0 300.915p 10000.0u 300.916p 0 301.115p 0 301.116p 10000.0u 301.117p 0 303.251p 0 303.252p 10000.0u 303.253p 0 309.662p 0 309.663p 10000.0u 309.664p 0 319.181p 0 319.182p 10000.0u 319.183p 0 320.147p 0 320.148p 10000.0u 320.149p 0 363.536p 0 363.537p 10000.0u 363.538p 0 364.454p 0 364.455p 10000.0u 364.456p 0 385.25p 0 385.251p 10000.0u 385.252p 0 399.092p 0 399.093p 10000.0u 399.094p 0 403.943p 0 403.944p 10000.0u 403.945p 0 411.86p 0 411.861p 10000.0u 411.862p 0 413.129p 0 413.13p 10000.0u 413.131p 0 414.353p 0 414.354p 10000.0u 414.355p 0 421.784p 0 421.785p 10000.0u 421.786p 0 434.288p 0 434.289p 10000.0u 434.29p 0 450.158p 0 450.159p 10000.0u 450.16p 0 472.367p 0 472.368p 10000.0u 472.369p 0 475.826p 0 475.827p 10000.0u 475.828p 0 480.809p 0 480.81p 10000.0u 480.811p 0 498.722p 0 498.723p 10000.0u 498.724p 0 499.442p 0 499.443p 10000.0u 499.444p 0 505.424p 0 505.425p 10000.0u 505.426p 0 512.129p 0 512.13p 10000.0u 512.131p 0 524.669p 0 524.67p 10000.0u 524.671p 0 528.29p 0 528.291p 10000.0u 528.292p 0 528.653p 0 528.654p 10000.0u 528.655p 0 558.872p 0 558.873p 10000.0u 558.874p 0 563.945p 0 563.946p 10000.0u 563.947p 0 565.076p 0 565.077p 10000.0u 565.078p 0 579.698p 0 579.699p 10000.0u 579.7p 0 582.764p 0 582.765p 10000.0u 582.766p 0 588.83p 0 588.831p 10000.0u 588.832p 0 608.189p 0 608.19p 10000.0u 608.191p 0 618.113p 0 618.114p 10000.0u 618.115p 0 620.183p 0 620.184p 10000.0u 620.185p 0 629.825p 0 629.826p 10000.0u 629.827p 0 631.508p 0 631.509p 10000.0u 631.51p 0 634.436p 0 634.437p 10000.0u 634.438p 0 643.649p 0 643.65p 10000.0u 643.651p 0 657.908p 0 657.909p 10000.0u 657.91p 0 658.658p 0 658.659p 10000.0u 658.66p 0 672.539p 0 672.54p 10000.0u 672.541p 0 676.283p 0 676.284p 10000.0u 676.285p 0 684.491p 0 684.492p 10000.0u 684.493p 0 693.557p 0 693.558p 10000.0u 693.559p 0 701.441p 0 701.442p 10000.0u 701.443p 0 704.897p 0 704.898p 10000.0u 704.899p 0 724.016p 0 724.017p 10000.0u 724.018p 0 731.225p 0 731.226p 10000.0u 731.227p 0 732.779p 0 732.78p 10000.0u 732.781p 0 750.566p 0 750.567p 10000.0u 750.568p 0 755.189p 0 755.19p 10000.0u 755.191p 0 756.074p 0 756.075p 10000.0u 756.076p 0 772.079p 0 772.08p 10000.0u 772.081p 0 774.818p 0 774.819p 10000.0u 774.82p 0 794.135p 0 794.136p 10000.0u 794.137p 0 802.214p 0 802.215p 10000.0u 802.216p 0 831.977p 0 831.978p 10000.0u 831.979p 0 834.068p 0 834.069p 10000.0u 834.07p 0 839.687p 0 839.688p 10000.0u 839.689p 0 867.785p 0 867.786p 10000.0u 867.787p 0 879.254p 0 879.255p 10000.0u 879.256p 0 885.272p 0 885.273p 10000.0u 885.274p 0 886.01p 0 886.011p 10000.0u 886.012p 0 892.355p 0 892.356p 10000.0u 892.357p 0 941.918p 0 941.919p 10000.0u 941.92p 0 943.589p 0 943.59p 10000.0u 943.591p 0 943.859p 0 943.86p 10000.0u 943.861p 0 955.649p 0 955.65p 10000.0u 955.651p 0 959.477p 0 959.478p 10000.0u 959.479p 0 969.236p 0 969.237p 10000.0u 969.238p 0 973.526p 0 973.527p 10000.0u 973.528p 0 982.664p 0 982.665p 10000.0u 982.666p 0 983.09p 0 983.091p 10000.0u 983.092p 0)
IIN63 0 64 pwl(0 0 24.965p 0 24.966p 10000.0u 24.967p 0 26.3p 0 26.301p 10000.0u 26.302p 0 52.823p 0 52.824p 10000.0u 52.825p 0 71.054p 0 71.055p 10000.0u 71.056p 0 82.028p 0 82.029p 10000.0u 82.03p 0 107.621p 0 107.622p 10000.0u 107.623p 0 114.842p 0 114.843p 10000.0u 114.844p 0 125.798p 0 125.799p 10000.0u 125.8p 0 133.676p 0 133.677p 10000.0u 133.678p 0 154.604p 0 154.605p 10000.0u 154.606p 0 158.588p 0 158.589p 10000.0u 158.59p 0 160.919p 0 160.92p 10000.0u 160.921p 0 166.412p 0 166.413p 10000.0u 166.414p 0 175.949p 0 175.95p 10000.0u 175.951p 0 190.592p 0 190.593p 10000.0u 190.594p 0 192.998p 0 192.999p 10000.0u 193.0p 0 200.219p 0 200.22p 10000.0u 200.221p 0 202.139p 0 202.14p 10000.0u 202.141p 0 237.509p 0 237.51p 10000.0u 237.511p 0 243.791p 0 243.792p 10000.0u 243.793p 0 248.726p 0 248.727p 10000.0u 248.728p 0 250.271p 0 250.272p 10000.0u 250.273p 0 251.822p 0 251.823p 10000.0u 251.824p 0 256.793p 0 256.794p 10000.0u 256.795p 0 270.419p 0 270.42p 10000.0u 270.421p 0 279.083p 0 279.084p 10000.0u 279.085p 0 286.409p 0 286.41p 10000.0u 286.411p 0 304.019p 0 304.02p 10000.0u 304.021p 0 305.444p 0 305.445p 10000.0u 305.446p 0 324.392p 0 324.393p 10000.0u 324.394p 0 327.44p 0 327.441p 10000.0u 327.442p 0 328.979p 0 328.98p 10000.0u 328.981p 0 329.999p 0 330.0p 10000.0u 330.001p 0 349.934p 0 349.935p 10000.0u 349.936p 0 356.834p 0 356.835p 10000.0u 356.836p 0 362.957p 0 362.958p 10000.0u 362.959p 0 365.192p 0 365.193p 10000.0u 365.194p 0 376.259p 0 376.26p 10000.0u 376.261p 0 387.683p 0 387.684p 10000.0u 387.685p 0 417.686p 0 417.687p 10000.0u 417.688p 0 424.16p 0 424.161p 10000.0u 424.162p 0 436.424p 0 436.425p 10000.0u 436.426p 0 437.546p 0 437.547p 10000.0u 437.548p 0 438.224p 0 438.225p 10000.0u 438.226p 0 452.156p 0 452.157p 10000.0u 452.158p 0 462.764p 0 462.765p 10000.0u 462.766p 0 471.758p 0 471.759p 10000.0u 471.76p 0 476.696p 0 476.697p 10000.0u 476.698p 0 491.102p 0 491.103p 10000.0u 491.104p 0 493.604p 0 493.605p 10000.0u 493.606p 0 493.874p 0 493.875p 10000.0u 493.876p 0 518.009p 0 518.01p 10000.0u 518.011p 0 529.679p 0 529.68p 10000.0u 529.681p 0 562.307p 0 562.308p 10000.0u 562.309p 0 564.305p 0 564.306p 10000.0u 564.307p 0 569.708p 0 569.709p 10000.0u 569.71p 0 570.56p 0 570.561p 10000.0u 570.562p 0 572.102p 0 572.103p 10000.0u 572.104p 0 572.75p 0 572.751p 10000.0u 572.752p 0 583.709p 0 583.71p 10000.0u 583.711p 0 610.574p 0 610.575p 10000.0u 610.576p 0 620.174p 0 620.175p 10000.0u 620.176p 0 635.291p 0 635.292p 10000.0u 635.293p 0 683.912p 0 683.913p 10000.0u 683.914p 0 697.202p 0 697.203p 10000.0u 697.204p 0 704.789p 0 704.79p 10000.0u 704.791p 0 715.775p 0 715.776p 10000.0u 715.777p 0 718.736p 0 718.737p 10000.0u 718.738p 0 735.071p 0 735.072p 10000.0u 735.073p 0 736.013p 0 736.014p 10000.0u 736.015p 0 747.263p 0 747.264p 10000.0u 747.265p 0 756.665p 0 756.666p 10000.0u 756.667p 0 760.565p 0 760.566p 10000.0u 760.567p 0 763.349p 0 763.35p 10000.0u 763.351p 0 764.453p 0 764.454p 10000.0u 764.455p 0 787.01p 0 787.011p 10000.0u 787.012p 0 789.23p 0 789.231p 10000.0u 789.232p 0 789.542p 0 789.543p 10000.0u 789.544p 0 790.754p 0 790.755p 10000.0u 790.756p 0 799.565p 0 799.566p 10000.0u 799.567p 0 807.623p 0 807.624p 10000.0u 807.625p 0 808.871p 0 808.872p 10000.0u 808.873p 0 811.574p 0 811.575p 10000.0u 811.576p 0 816.503p 0 816.504p 10000.0u 816.505p 0 823.304p 0 823.305p 10000.0u 823.306p 0 847.817p 0 847.818p 10000.0u 847.819p 0 856.103p 0 856.104p 10000.0u 856.105p 0 863.003p 0 863.004p 10000.0u 863.005p 0 863.732p 0 863.733p 10000.0u 863.734p 0 872.012p 0 872.013p 10000.0u 872.014p 0 872.588p 0 872.589p 10000.0u 872.59p 0 915.278p 0 915.279p 10000.0u 915.28p 0 920.591p 0 920.592p 10000.0u 920.593p 0 924.353p 0 924.354p 10000.0u 924.355p 0 937.589p 0 937.59p 10000.0u 937.591p 0 940.274p 0 940.275p 10000.0u 940.276p 0 947.714p 0 947.715p 10000.0u 947.716p 0 947.885p 0 947.886p 10000.0u 947.887p 0 948.839p 0 948.84p 10000.0u 948.841p 0 954.602p 0 954.603p 10000.0u 954.604p 0 961.772p 0 961.773p 10000.0u 961.774p 0 974.327p 0 974.328p 10000.0u 974.329p 0 974.612p 0 974.613p 10000.0u 974.614p 0 978.452p 0 978.453p 10000.0u 978.454p 0 979.283p 0 979.284p 10000.0u 979.285p 0 982.919p 0 982.92p 10000.0u 982.921p 0)
IIN64 0 65 pwl(0 0 18.98p 0 18.981p 10000.0u 18.982p 0 46.769p 0 46.77p 10000.0u 46.771p 0 60.14p 0 60.141p 10000.0u 60.142p 0 62.996p 0 62.997p 10000.0u 62.998p 0 64.991p 0 64.992p 10000.0u 64.993p 0 71.651p 0 71.652p 10000.0u 71.653p 0 99.407p 0 99.408p 10000.0u 99.409p 0 113.345p 0 113.346p 10000.0u 113.347p 0 117.335p 0 117.336p 10000.0u 117.337p 0 128.093p 0 128.094p 10000.0u 128.095p 0 140.981p 0 140.982p 10000.0u 140.983p 0 141.704p 0 141.705p 10000.0u 141.706p 0 144.626p 0 144.627p 10000.0u 144.628p 0 153.641p 0 153.642p 10000.0u 153.643p 0 192.5p 0 192.501p 10000.0u 192.502p 0 207.425p 0 207.426p 10000.0u 207.427p 0 211.508p 0 211.509p 10000.0u 211.51p 0 211.586p 0 211.587p 10000.0u 211.588p 0 222.485p 0 222.486p 10000.0u 222.487p 0 225.659p 0 225.66p 10000.0u 225.661p 0 264.467p 0 264.468p 10000.0u 264.469p 0 270.368p 0 270.369p 10000.0u 270.37p 0 300.359p 0 300.36p 10000.0u 300.361p 0 306.749p 0 306.75p 10000.0u 306.751p 0 312.659p 0 312.66p 10000.0u 312.661p 0 325.88p 0 325.881p 10000.0u 325.882p 0 328.457p 0 328.458p 10000.0u 328.459p 0 337.403p 0 337.404p 10000.0u 337.405p 0 385.784p 0 385.785p 10000.0u 385.786p 0 396.188p 0 396.189p 10000.0u 396.19p 0 406.499p 0 406.5p 10000.0u 406.501p 0 411.407p 0 411.408p 10000.0u 411.409p 0 416.879p 0 416.88p 10000.0u 416.881p 0 448.904p 0 448.905p 10000.0u 448.906p 0 451.643p 0 451.644p 10000.0u 451.645p 0 482.987p 0 482.988p 10000.0u 482.989p 0 505.694p 0 505.695p 10000.0u 505.696p 0 511.613p 0 511.614p 10000.0u 511.615p 0 518.126p 0 518.127p 10000.0u 518.128p 0 519.557p 0 519.558p 10000.0u 519.559p 0 520.547p 0 520.548p 10000.0u 520.549p 0 532.505p 0 532.506p 10000.0u 532.507p 0 549.959p 0 549.96p 10000.0u 549.961p 0 555.296p 0 555.297p 10000.0u 555.298p 0 567.341p 0 567.342p 10000.0u 567.343p 0 585.581p 0 585.582p 10000.0u 585.583p 0 603.167p 0 603.168p 10000.0u 603.169p 0 617.486p 0 617.487p 10000.0u 617.488p 0 623.669p 0 623.67p 10000.0u 623.671p 0 639.599p 0 639.6p 10000.0u 639.601p 0 643.307p 0 643.308p 10000.0u 643.309p 0 648.29p 0 648.291p 10000.0u 648.292p 0 661.562p 0 661.563p 10000.0u 661.564p 0 665.09p 0 665.091p 10000.0u 665.092p 0 683.732p 0 683.733p 10000.0u 683.734p 0 685.754p 0 685.755p 10000.0u 685.756p 0 695.396p 0 695.397p 10000.0u 695.398p 0 726.485p 0 726.486p 10000.0u 726.487p 0 727.622p 0 727.623p 10000.0u 727.624p 0 742.568p 0 742.569p 10000.0u 742.57p 0 758.072p 0 758.073p 10000.0u 758.074p 0 761.495p 0 761.496p 10000.0u 761.497p 0 763.619p 0 763.62p 10000.0u 763.621p 0 768.212p 0 768.213p 10000.0u 768.214p 0 781.748p 0 781.749p 10000.0u 781.75p 0 790.766p 0 790.767p 10000.0u 790.768p 0 801.134p 0 801.135p 10000.0u 801.136p 0 803.462p 0 803.463p 10000.0u 803.464p 0 811.31p 0 811.311p 10000.0u 811.312p 0 815.747p 0 815.748p 10000.0u 815.749p 0 831.314p 0 831.315p 10000.0u 831.316p 0 833.432p 0 833.433p 10000.0u 833.434p 0 837.314p 0 837.315p 10000.0u 837.316p 0 848.36p 0 848.361p 10000.0u 848.362p 0 851.105p 0 851.106p 10000.0u 851.107p 0 851.324p 0 851.325p 10000.0u 851.326p 0 855.968p 0 855.969p 10000.0u 855.97p 0 875.828p 0 875.829p 10000.0u 875.83p 0 897.617p 0 897.618p 10000.0u 897.619p 0 906.326p 0 906.327p 10000.0u 906.328p 0 908.162p 0 908.163p 10000.0u 908.164p 0 925.07p 0 925.071p 10000.0u 925.072p 0 928.859p 0 928.86p 10000.0u 928.861p 0 936.803p 0 936.804p 10000.0u 936.805p 0 942.695p 0 942.696p 10000.0u 942.697p 0 951.434p 0 951.435p 10000.0u 951.436p 0 956.195p 0 956.196p 10000.0u 956.197p 0 959.57p 0 959.571p 10000.0u 959.572p 0 979.277p 0 979.278p 10000.0u 979.279p 0 998.579p 0 998.58p 10000.0u 998.581p 0)
IIN65 0 66 pwl(0 0 2.708p 0 2.709p 10000.0u 2.71p 0 10.217p 0 10.218p 10000.0u 10.219p 0 25.364p 0 25.365p 10000.0u 25.366p 0 29.966p 0 29.967p 10000.0u 29.968p 0 37.22p 0 37.221p 10000.0u 37.222p 0 40.835p 0 40.836p 10000.0u 40.837p 0 51.635p 0 51.636p 10000.0u 51.637p 0 63.224p 0 63.225p 10000.0u 63.226p 0 66.671p 0 66.672p 10000.0u 66.673p 0 100.679p 0 100.68p 10000.0u 100.681p 0 122.903p 0 122.904p 10000.0u 122.905p 0 124.859p 0 124.86p 10000.0u 124.861p 0 140.945p 0 140.946p 10000.0u 140.947p 0 154.037p 0 154.038p 10000.0u 154.039p 0 156.32p 0 156.321p 10000.0u 156.322p 0 163.469p 0 163.47p 10000.0u 163.471p 0 164.945p 0 164.946p 10000.0u 164.947p 0 165.908p 0 165.909p 10000.0u 165.91p 0 175.184p 0 175.185p 10000.0u 175.186p 0 185.9p 0 185.901p 10000.0u 185.902p 0 188.768p 0 188.769p 10000.0u 188.77p 0 195.68p 0 195.681p 10000.0u 195.682p 0 203.954p 0 203.955p 10000.0u 203.956p 0 211.049p 0 211.05p 10000.0u 211.051p 0 213.233p 0 213.234p 10000.0u 213.235p 0 234.395p 0 234.396p 10000.0u 234.397p 0 238.88p 0 238.881p 10000.0u 238.882p 0 252.596p 0 252.597p 10000.0u 252.598p 0 254.066p 0 254.067p 10000.0u 254.068p 0 254.183p 0 254.184p 10000.0u 254.185p 0 277.706p 0 277.707p 10000.0u 277.708p 0 280.184p 0 280.185p 10000.0u 280.186p 0 293.807p 0 293.808p 10000.0u 293.809p 0 297.08p 0 297.081p 10000.0u 297.082p 0 301.94p 0 301.941p 10000.0u 301.942p 0 302.984p 0 302.985p 10000.0u 302.986p 0 318.08p 0 318.081p 10000.0u 318.082p 0 345.461p 0 345.462p 10000.0u 345.463p 0 369.56p 0 369.561p 10000.0u 369.562p 0 390.971p 0 390.972p 10000.0u 390.973p 0 398.765p 0 398.766p 10000.0u 398.767p 0 404.48p 0 404.481p 10000.0u 404.482p 0 405.329p 0 405.33p 10000.0u 405.331p 0 407.288p 0 407.289p 10000.0u 407.29p 0 410.168p 0 410.169p 10000.0u 410.17p 0 431.816p 0 431.817p 10000.0u 431.818p 0 433.331p 0 433.332p 10000.0u 433.333p 0 465.584p 0 465.585p 10000.0u 465.586p 0 468.77p 0 468.771p 10000.0u 468.772p 0 474.719p 0 474.72p 10000.0u 474.721p 0 475.637p 0 475.638p 10000.0u 475.639p 0 488.204p 0 488.205p 10000.0u 488.206p 0 490.604p 0 490.605p 10000.0u 490.606p 0 499.43p 0 499.431p 10000.0u 499.432p 0 507.155p 0 507.156p 10000.0u 507.157p 0 519.08p 0 519.081p 10000.0u 519.082p 0 539.324p 0 539.325p 10000.0u 539.326p 0 566.066p 0 566.067p 10000.0u 566.068p 0 585.38p 0 585.381p 10000.0u 585.382p 0 585.542p 0 585.543p 10000.0u 585.544p 0 587.015p 0 587.016p 10000.0u 587.017p 0 592.217p 0 592.218p 10000.0u 592.219p 0 597.923p 0 597.924p 10000.0u 597.925p 0 609.044p 0 609.045p 10000.0u 609.046p 0 621.08p 0 621.081p 10000.0u 621.082p 0 621.611p 0 621.612p 10000.0u 621.613p 0 621.842p 0 621.843p 10000.0u 621.844p 0 624.095p 0 624.096p 10000.0u 624.097p 0 640.016p 0 640.017p 10000.0u 640.018p 0 649.547p 0 649.548p 10000.0u 649.549p 0 662.303p 0 662.304p 10000.0u 662.305p 0 664.196p 0 664.197p 10000.0u 664.198p 0 666.392p 0 666.393p 10000.0u 666.394p 0 694.997p 0 694.998p 10000.0u 694.999p 0 718.979p 0 718.98p 10000.0u 718.981p 0 724.013p 0 724.014p 10000.0u 724.015p 0 752.312p 0 752.313p 10000.0u 752.314p 0 771.188p 0 771.189p 10000.0u 771.19p 0 795.335p 0 795.336p 10000.0u 795.337p 0 797.705p 0 797.706p 10000.0u 797.707p 0 800.105p 0 800.106p 10000.0u 800.107p 0 829.979p 0 829.98p 10000.0u 829.981p 0 836.537p 0 836.538p 10000.0u 836.539p 0 844.535p 0 844.536p 10000.0u 844.537p 0 859.127p 0 859.128p 10000.0u 859.129p 0 862.409p 0 862.41p 10000.0u 862.411p 0 868.508p 0 868.509p 10000.0u 868.51p 0 874.967p 0 874.968p 10000.0u 874.969p 0 877.559p 0 877.56p 10000.0u 877.561p 0 882.536p 0 882.537p 10000.0u 882.538p 0 888.824p 0 888.825p 10000.0u 888.826p 0 898.661p 0 898.662p 10000.0u 898.663p 0 913.715p 0 913.716p 10000.0u 913.717p 0 914.546p 0 914.547p 10000.0u 914.548p 0 939.809p 0 939.81p 10000.0u 939.811p 0 943.913p 0 943.914p 10000.0u 943.915p 0 990.329p 0 990.33p 10000.0u 990.331p 0 992.345p 0 992.346p 10000.0u 992.347p 0 993.401p 0 993.402p 10000.0u 993.403p 0)
IIN66 0 67 pwl(0 0 0.566p 0 0.567p 10000.0u 0.568p 0 4.205p 0 4.206p 10000.0u 4.207p 0 7.508p 0 7.509p 10000.0u 7.51p 0 13.361p 0 13.362p 10000.0u 13.363p 0 32.459p 0 32.46p 10000.0u 32.461p 0 47.9p 0 47.901p 10000.0u 47.902p 0 49.217p 0 49.218p 10000.0u 49.219p 0 108.863p 0 108.864p 10000.0u 108.865p 0 114.188p 0 114.189p 10000.0u 114.19p 0 122.006p 0 122.007p 10000.0u 122.008p 0 140.825p 0 140.826p 10000.0u 140.827p 0 158.081p 0 158.082p 10000.0u 158.083p 0 162.935p 0 162.936p 10000.0u 162.937p 0 175.949p 0 175.95p 10000.0u 175.951p 0 198.038p 0 198.039p 10000.0u 198.04p 0 199.337p 0 199.338p 10000.0u 199.339p 0 201.455p 0 201.456p 10000.0u 201.457p 0 202.718p 0 202.719p 10000.0u 202.72p 0 205.193p 0 205.194p 10000.0u 205.195p 0 216.266p 0 216.267p 10000.0u 216.268p 0 234.098p 0 234.099p 10000.0u 234.1p 0 235.307p 0 235.308p 10000.0u 235.309p 0 240.218p 0 240.219p 10000.0u 240.22p 0 246.482p 0 246.483p 10000.0u 246.484p 0 250.655p 0 250.656p 10000.0u 250.657p 0 252.323p 0 252.324p 10000.0u 252.325p 0 253.532p 0 253.533p 10000.0u 253.534p 0 269.786p 0 269.787p 10000.0u 269.788p 0 272.168p 0 272.169p 10000.0u 272.17p 0 294.344p 0 294.345p 10000.0u 294.346p 0 314.186p 0 314.187p 10000.0u 314.188p 0 326.252p 0 326.253p 10000.0u 326.254p 0 344.801p 0 344.802p 10000.0u 344.803p 0 360.842p 0 360.843p 10000.0u 360.844p 0 385.355p 0 385.356p 10000.0u 385.357p 0 393.44p 0 393.441p 10000.0u 393.442p 0 421.547p 0 421.548p 10000.0u 421.549p 0 425.048p 0 425.049p 10000.0u 425.05p 0 427.025p 0 427.026p 10000.0u 427.027p 0 433.07p 0 433.071p 10000.0u 433.072p 0 443.591p 0 443.592p 10000.0u 443.593p 0 444.428p 0 444.429p 10000.0u 444.43p 0 455.411p 0 455.412p 10000.0u 455.413p 0 463.718p 0 463.719p 10000.0u 463.72p 0 467.354p 0 467.355p 10000.0u 467.356p 0 472.238p 0 472.239p 10000.0u 472.24p 0 475.202p 0 475.203p 10000.0u 475.204p 0 490.997p 0 490.998p 10000.0u 490.999p 0 503.945p 0 503.946p 10000.0u 503.947p 0 507.725p 0 507.726p 10000.0u 507.727p 0 510.284p 0 510.285p 10000.0u 510.286p 0 522.188p 0 522.189p 10000.0u 522.19p 0 534.248p 0 534.249p 10000.0u 534.25p 0 545.978p 0 545.979p 10000.0u 545.98p 0 566.855p 0 566.856p 10000.0u 566.857p 0 568.682p 0 568.683p 10000.0u 568.684p 0 569.0p 0 569.001p 10000.0u 569.002p 0 594.605p 0 594.606p 10000.0u 594.607p 0 594.998p 0 594.999p 10000.0u 595.0p 0 607.718p 0 607.719p 10000.0u 607.72p 0 611.213p 0 611.214p 10000.0u 611.215p 0 622.739p 0 622.74p 10000.0u 622.741p 0 625.682p 0 625.683p 10000.0u 625.684p 0 627.62p 0 627.621p 10000.0u 627.622p 0 644.75p 0 644.751p 10000.0u 644.752p 0 650.051p 0 650.052p 10000.0u 650.053p 0 655.403p 0 655.404p 10000.0u 655.405p 0 657.341p 0 657.342p 10000.0u 657.343p 0 670.466p 0 670.467p 10000.0u 670.468p 0 680.06p 0 680.061p 10000.0u 680.062p 0 691.718p 0 691.719p 10000.0u 691.72p 0 698.558p 0 698.559p 10000.0u 698.56p 0 734.375p 0 734.376p 10000.0u 734.377p 0 747.212p 0 747.213p 10000.0u 747.214p 0 751.352p 0 751.353p 10000.0u 751.354p 0 751.886p 0 751.887p 10000.0u 751.888p 0 755.549p 0 755.55p 10000.0u 755.551p 0 756.086p 0 756.087p 10000.0u 756.088p 0 765.689p 0 765.69p 10000.0u 765.691p 0 769.877p 0 769.878p 10000.0u 769.879p 0 784.61p 0 784.611p 10000.0u 784.612p 0 788.597p 0 788.598p 10000.0u 788.599p 0 799.34p 0 799.341p 10000.0u 799.342p 0 802.457p 0 802.458p 10000.0u 802.459p 0 818.063p 0 818.064p 10000.0u 818.065p 0 839.444p 0 839.445p 10000.0u 839.446p 0 849.449p 0 849.45p 10000.0u 849.451p 0 873.032p 0 873.033p 10000.0u 873.034p 0 873.425p 0 873.426p 10000.0u 873.427p 0 877.076p 0 877.077p 10000.0u 877.078p 0 891.341p 0 891.342p 10000.0u 891.343p 0 891.716p 0 891.717p 10000.0u 891.718p 0 902.558p 0 902.559p 10000.0u 902.56p 0 923.309p 0 923.31p 10000.0u 923.311p 0 932.489p 0 932.49p 10000.0u 932.491p 0 950.684p 0 950.685p 10000.0u 950.686p 0 957.911p 0 957.912p 10000.0u 957.913p 0 961.67p 0 961.671p 10000.0u 961.672p 0 978.488p 0 978.489p 10000.0u 978.49p 0 978.839p 0 978.84p 10000.0u 978.841p 0 982.487p 0 982.488p 10000.0u 982.489p 0)
IIN67 0 68 pwl(0 0 56.726p 0 56.727p 10000.0u 56.728p 0 69.833p 0 69.834p 10000.0u 69.835p 0 132.917p 0 132.918p 10000.0u 132.919p 0 133.4p 0 133.401p 10000.0u 133.402p 0 136.721p 0 136.722p 10000.0u 136.723p 0 140.387p 0 140.388p 10000.0u 140.389p 0 142.433p 0 142.434p 10000.0u 142.435p 0 142.91p 0 142.911p 10000.0u 142.912p 0 143.114p 0 143.115p 10000.0u 143.116p 0 144.611p 0 144.612p 10000.0u 144.613p 0 158.729p 0 158.73p 10000.0u 158.731p 0 160.106p 0 160.107p 10000.0u 160.108p 0 164.75p 0 164.751p 10000.0u 164.752p 0 168.101p 0 168.102p 10000.0u 168.103p 0 169.196p 0 169.197p 10000.0u 169.198p 0 202.616p 0 202.617p 10000.0u 202.618p 0 206.183p 0 206.184p 10000.0u 206.185p 0 213.047p 0 213.048p 10000.0u 213.049p 0 230.888p 0 230.889p 10000.0u 230.89p 0 246.011p 0 246.012p 10000.0u 246.013p 0 261.314p 0 261.315p 10000.0u 261.316p 0 263.375p 0 263.376p 10000.0u 263.377p 0 264.524p 0 264.525p 10000.0u 264.526p 0 266.813p 0 266.814p 10000.0u 266.815p 0 276.575p 0 276.576p 10000.0u 276.577p 0 282.416p 0 282.417p 10000.0u 282.418p 0 287.66p 0 287.661p 10000.0u 287.662p 0 292.163p 0 292.164p 10000.0u 292.165p 0 303.794p 0 303.795p 10000.0u 303.796p 0 307.103p 0 307.104p 10000.0u 307.105p 0 315.476p 0 315.477p 10000.0u 315.478p 0 321.347p 0 321.348p 10000.0u 321.349p 0 322.517p 0 322.518p 10000.0u 322.519p 0 325.844p 0 325.845p 10000.0u 325.846p 0 329.546p 0 329.547p 10000.0u 329.548p 0 333.635p 0 333.636p 10000.0u 333.637p 0 356.147p 0 356.148p 10000.0u 356.149p 0 356.222p 0 356.223p 10000.0u 356.224p 0 361.565p 0 361.566p 10000.0u 361.567p 0 377.774p 0 377.775p 10000.0u 377.776p 0 381.515p 0 381.516p 10000.0u 381.517p 0 402.32p 0 402.321p 10000.0u 402.322p 0 404.663p 0 404.664p 10000.0u 404.665p 0 407.924p 0 407.925p 10000.0u 407.926p 0 417.413p 0 417.414p 10000.0u 417.415p 0 422.096p 0 422.097p 10000.0u 422.098p 0 454.163p 0 454.164p 10000.0u 454.165p 0 483.851p 0 483.852p 10000.0u 483.853p 0 483.86p 0 483.861p 10000.0u 483.862p 0 513.665p 0 513.666p 10000.0u 513.667p 0 518.642p 0 518.643p 10000.0u 518.644p 0 523.634p 0 523.635p 10000.0u 523.636p 0 539.861p 0 539.862p 10000.0u 539.863p 0 549.776p 0 549.777p 10000.0u 549.778p 0 553.895p 0 553.896p 10000.0u 553.897p 0 557.237p 0 557.238p 10000.0u 557.239p 0 565.583p 0 565.584p 10000.0u 565.585p 0 579.092p 0 579.093p 10000.0u 579.094p 0 579.254p 0 579.255p 10000.0u 579.256p 0 601.694p 0 601.695p 10000.0u 601.696p 0 603.428p 0 603.429p 10000.0u 603.43p 0 615.023p 0 615.024p 10000.0u 615.025p 0 629.783p 0 629.784p 10000.0u 629.785p 0 639.485p 0 639.486p 10000.0u 639.487p 0 641.96p 0 641.961p 10000.0u 641.962p 0 643.331p 0 643.332p 10000.0u 643.333p 0 658.826p 0 658.827p 10000.0u 658.828p 0 662.099p 0 662.1p 10000.0u 662.101p 0 663.458p 0 663.459p 10000.0u 663.46p 0 665.036p 0 665.037p 10000.0u 665.038p 0 666.413p 0 666.414p 10000.0u 666.415p 0 685.22p 0 685.221p 10000.0u 685.222p 0 688.286p 0 688.287p 10000.0u 688.288p 0 694.439p 0 694.44p 10000.0u 694.441p 0 697.805p 0 697.806p 10000.0u 697.807p 0 699.194p 0 699.195p 10000.0u 699.196p 0 699.806p 0 699.807p 10000.0u 699.808p 0 704.993p 0 704.994p 10000.0u 704.995p 0 719.27p 0 719.271p 10000.0u 719.272p 0 735.899p 0 735.9p 10000.0u 735.901p 0 740.837p 0 740.838p 10000.0u 740.839p 0 758.411p 0 758.412p 10000.0u 758.413p 0 759.122p 0 759.123p 10000.0u 759.124p 0 769.619p 0 769.62p 10000.0u 769.621p 0 780.692p 0 780.693p 10000.0u 780.694p 0 781.235p 0 781.236p 10000.0u 781.237p 0 782.333p 0 782.334p 10000.0u 782.335p 0 783.746p 0 783.747p 10000.0u 783.748p 0 793.118p 0 793.119p 10000.0u 793.12p 0 794.414p 0 794.415p 10000.0u 794.416p 0 799.604p 0 799.605p 10000.0u 799.606p 0 817.484p 0 817.485p 10000.0u 817.486p 0 835.994p 0 835.995p 10000.0u 835.996p 0 856.718p 0 856.719p 10000.0u 856.72p 0 897.245p 0 897.246p 10000.0u 897.247p 0 903.299p 0 903.3p 10000.0u 903.301p 0 908.861p 0 908.862p 10000.0u 908.863p 0 912.731p 0 912.732p 10000.0u 912.733p 0 913.169p 0 913.17p 10000.0u 913.171p 0 927.998p 0 927.999p 10000.0u 928.0p 0 930.131p 0 930.132p 10000.0u 930.133p 0 944.576p 0 944.577p 10000.0u 944.578p 0 960.734p 0 960.735p 10000.0u 960.736p 0 970.178p 0 970.179p 10000.0u 970.18p 0 975.017p 0 975.018p 10000.0u 975.019p 0 978.29p 0 978.291p 10000.0u 978.292p 0 991.688p 0 991.689p 10000.0u 991.69p 0)
IIN68 0 69 pwl(0 0 0.047p 0 0.048p 10000.0u 0.049p 0 3.269p 0 3.27p 10000.0u 3.271p 0 13.607p 0 13.608p 10000.0u 13.609p 0 18.563p 0 18.564p 10000.0u 18.565p 0 30.137p 0 30.138p 10000.0u 30.139p 0 40.715p 0 40.716p 10000.0u 40.717p 0 41.684p 0 41.685p 10000.0u 41.686p 0 62.696p 0 62.697p 10000.0u 62.698p 0 69.389p 0 69.39p 10000.0u 69.391p 0 73.364p 0 73.365p 10000.0u 73.366p 0 89.456p 0 89.457p 10000.0u 89.458p 0 90.581p 0 90.582p 10000.0u 90.583p 0 114.944p 0 114.945p 10000.0u 114.946p 0 124.772p 0 124.773p 10000.0u 124.774p 0 132.578p 0 132.579p 10000.0u 132.58p 0 133.034p 0 133.035p 10000.0u 133.036p 0 135.602p 0 135.603p 10000.0u 135.604p 0 146.519p 0 146.52p 10000.0u 146.521p 0 174.131p 0 174.132p 10000.0u 174.133p 0 190.922p 0 190.923p 10000.0u 190.924p 0 206.642p 0 206.643p 10000.0u 206.644p 0 207.413p 0 207.414p 10000.0u 207.415p 0 212.267p 0 212.268p 10000.0u 212.269p 0 215.906p 0 215.907p 10000.0u 215.908p 0 217.079p 0 217.08p 10000.0u 217.081p 0 225.278p 0 225.279p 10000.0u 225.28p 0 230.132p 0 230.133p 10000.0u 230.134p 0 236.687p 0 236.688p 10000.0u 236.689p 0 244.787p 0 244.788p 10000.0u 244.789p 0 252.257p 0 252.258p 10000.0u 252.259p 0 256.058p 0 256.059p 10000.0u 256.06p 0 260.288p 0 260.289p 10000.0u 260.29p 0 262.559p 0 262.56p 10000.0u 262.561p 0 271.082p 0 271.083p 10000.0u 271.084p 0 275.108p 0 275.109p 10000.0u 275.11p 0 275.645p 0 275.646p 10000.0u 275.647p 0 284.945p 0 284.946p 10000.0u 284.947p 0 285.467p 0 285.468p 10000.0u 285.469p 0 290.054p 0 290.055p 10000.0u 290.056p 0 293.636p 0 293.637p 10000.0u 293.638p 0 295.577p 0 295.578p 10000.0u 295.579p 0 341.222p 0 341.223p 10000.0u 341.224p 0 345.161p 0 345.162p 10000.0u 345.163p 0 349.277p 0 349.278p 10000.0u 349.279p 0 354.497p 0 354.498p 10000.0u 354.499p 0 404.426p 0 404.427p 10000.0u 404.428p 0 405.221p 0 405.222p 10000.0u 405.223p 0 412.919p 0 412.92p 10000.0u 412.921p 0 425.417p 0 425.418p 10000.0u 425.419p 0 429.527p 0 429.528p 10000.0u 429.529p 0 437.108p 0 437.109p 10000.0u 437.11p 0 438.224p 0 438.225p 10000.0u 438.226p 0 438.863p 0 438.864p 10000.0u 438.865p 0 442.733p 0 442.734p 10000.0u 442.735p 0 445.826p 0 445.827p 10000.0u 445.828p 0 473.618p 0 473.619p 10000.0u 473.62p 0 517.715p 0 517.716p 10000.0u 517.717p 0 530.633p 0 530.634p 10000.0u 530.635p 0 541.256p 0 541.257p 10000.0u 541.258p 0 587.786p 0 587.787p 10000.0u 587.788p 0 612.191p 0 612.192p 10000.0u 612.193p 0 614.399p 0 614.4p 10000.0u 614.401p 0 618.74p 0 618.741p 10000.0u 618.742p 0 621.041p 0 621.042p 10000.0u 621.043p 0 621.833p 0 621.834p 10000.0u 621.835p 0 634.208p 0 634.209p 10000.0u 634.21p 0 635.363p 0 635.364p 10000.0u 635.365p 0 645.899p 0 645.9p 10000.0u 645.901p 0 668.09p 0 668.091p 10000.0u 668.092p 0 672.014p 0 672.015p 10000.0u 672.016p 0 706.157p 0 706.158p 10000.0u 706.159p 0 721.709p 0 721.71p 10000.0u 721.711p 0 729.359p 0 729.36p 10000.0u 729.361p 0 742.616p 0 742.617p 10000.0u 742.618p 0 769.16p 0 769.161p 10000.0u 769.162p 0 771.335p 0 771.336p 10000.0u 771.337p 0 792.68p 0 792.681p 10000.0u 792.682p 0 798.098p 0 798.099p 10000.0u 798.1p 0 819.668p 0 819.669p 10000.0u 819.67p 0 820.073p 0 820.074p 10000.0u 820.075p 0 825.443p 0 825.444p 10000.0u 825.445p 0 831.824p 0 831.825p 10000.0u 831.826p 0 835.529p 0 835.53p 10000.0u 835.531p 0 845.93p 0 845.931p 10000.0u 845.932p 0 849.692p 0 849.693p 10000.0u 849.694p 0 874.175p 0 874.176p 10000.0u 874.177p 0 876.257p 0 876.258p 10000.0u 876.259p 0 895.919p 0 895.92p 10000.0u 895.921p 0 908.072p 0 908.073p 10000.0u 908.074p 0 914.162p 0 914.163p 10000.0u 914.164p 0 936.092p 0 936.093p 10000.0u 936.094p 0 961.37p 0 961.371p 10000.0u 961.372p 0 965.732p 0 965.733p 10000.0u 965.734p 0 966.194p 0 966.195p 10000.0u 966.196p 0 969.002p 0 969.003p 10000.0u 969.004p 0 980.105p 0 980.106p 10000.0u 980.107p 0 980.255p 0 980.256p 10000.0u 980.257p 0 983.756p 0 983.757p 10000.0u 983.758p 0 998.765p 0 998.766p 10000.0u 998.767p 0)
IIN69 0 70 pwl(0 0 3.275p 0 3.276p 10000.0u 3.277p 0 7.07p 0 7.071p 10000.0u 7.072p 0 10.802p 0 10.803p 10000.0u 10.804p 0 10.988p 0 10.989p 10000.0u 10.99p 0 21.857p 0 21.858p 10000.0u 21.859p 0 49.469p 0 49.47p 10000.0u 49.471p 0 56.816p 0 56.817p 10000.0u 56.818p 0 70.496p 0 70.497p 10000.0u 70.498p 0 71.42p 0 71.421p 10000.0u 71.422p 0 93.593p 0 93.594p 10000.0u 93.595p 0 96.272p 0 96.273p 10000.0u 96.274p 0 98.675p 0 98.676p 10000.0u 98.677p 0 98.816p 0 98.817p 10000.0u 98.818p 0 113.114p 0 113.115p 10000.0u 113.116p 0 127.958p 0 127.959p 10000.0u 127.96p 0 131.156p 0 131.157p 10000.0u 131.158p 0 155.453p 0 155.454p 10000.0u 155.455p 0 179.885p 0 179.886p 10000.0u 179.887p 0 182.072p 0 182.073p 10000.0u 182.074p 0 187.136p 0 187.137p 10000.0u 187.138p 0 204.125p 0 204.126p 10000.0u 204.127p 0 212.192p 0 212.193p 10000.0u 212.194p 0 212.408p 0 212.409p 10000.0u 212.41p 0 239.567p 0 239.568p 10000.0u 239.569p 0 240.164p 0 240.165p 10000.0u 240.166p 0 243.083p 0 243.084p 10000.0u 243.085p 0 249.506p 0 249.507p 10000.0u 249.508p 0 261.782p 0 261.783p 10000.0u 261.784p 0 266.843p 0 266.844p 10000.0u 266.845p 0 277.652p 0 277.653p 10000.0u 277.654p 0 282.671p 0 282.672p 10000.0u 282.673p 0 294.152p 0 294.153p 10000.0u 294.154p 0 300.887p 0 300.888p 10000.0u 300.889p 0 307.304p 0 307.305p 10000.0u 307.306p 0 313.061p 0 313.062p 10000.0u 313.063p 0 327.554p 0 327.555p 10000.0u 327.556p 0 346.586p 0 346.587p 10000.0u 346.588p 0 368.165p 0 368.166p 10000.0u 368.167p 0 369.605p 0 369.606p 10000.0u 369.607p 0 379.022p 0 379.023p 10000.0u 379.024p 0 386.759p 0 386.76p 10000.0u 386.761p 0 407.558p 0 407.559p 10000.0u 407.56p 0 410.27p 0 410.271p 10000.0u 410.272p 0 417.299p 0 417.3p 10000.0u 417.301p 0 421.541p 0 421.542p 10000.0u 421.543p 0 426.563p 0 426.564p 10000.0u 426.565p 0 430.538p 0 430.539p 10000.0u 430.54p 0 440.168p 0 440.169p 10000.0u 440.17p 0 442.961p 0 442.962p 10000.0u 442.963p 0 446.558p 0 446.559p 10000.0u 446.56p 0 462.302p 0 462.303p 10000.0u 462.304p 0 472.592p 0 472.593p 10000.0u 472.594p 0 480.785p 0 480.786p 10000.0u 480.787p 0 493.355p 0 493.356p 10000.0u 493.357p 0 505.187p 0 505.188p 10000.0u 505.189p 0 505.502p 0 505.503p 10000.0u 505.504p 0 536.762p 0 536.763p 10000.0u 536.764p 0 537.434p 0 537.435p 10000.0u 537.436p 0 540.806p 0 540.807p 10000.0u 540.808p 0 541.997p 0 541.998p 10000.0u 541.999p 0 558.134p 0 558.135p 10000.0u 558.136p 0 559.229p 0 559.23p 10000.0u 559.231p 0 573.47p 0 573.471p 10000.0u 573.472p 0 575.513p 0 575.514p 10000.0u 575.515p 0 587.867p 0 587.868p 10000.0u 587.869p 0 592.262p 0 592.263p 10000.0u 592.264p 0 596.57p 0 596.571p 10000.0u 596.572p 0 599.399p 0 599.4p 10000.0u 599.401p 0 600.152p 0 600.153p 10000.0u 600.154p 0 609.38p 0 609.381p 10000.0u 609.382p 0 617.18p 0 617.181p 10000.0u 617.182p 0 632.621p 0 632.622p 10000.0u 632.623p 0 637.472p 0 637.473p 10000.0u 637.474p 0 638.066p 0 638.067p 10000.0u 638.068p 0 638.102p 0 638.103p 10000.0u 638.104p 0 642.572p 0 642.573p 10000.0u 642.574p 0 656.822p 0 656.823p 10000.0u 656.824p 0 675.311p 0 675.312p 10000.0u 675.313p 0 682.634p 0 682.635p 10000.0u 682.636p 0 684.335p 0 684.336p 10000.0u 684.337p 0 699.113p 0 699.114p 10000.0u 699.115p 0 737.69p 0 737.691p 10000.0u 737.692p 0 747.551p 0 747.552p 10000.0u 747.553p 0 748.928p 0 748.929p 10000.0u 748.93p 0 749.069p 0 749.07p 10000.0u 749.071p 0 751.907p 0 751.908p 10000.0u 751.909p 0 777.083p 0 777.084p 10000.0u 777.085p 0 789.323p 0 789.324p 10000.0u 789.325p 0 830.522p 0 830.523p 10000.0u 830.524p 0 833.405p 0 833.406p 10000.0u 833.407p 0 841.154p 0 841.155p 10000.0u 841.156p 0 847.283p 0 847.284p 10000.0u 847.285p 0 860.345p 0 860.346p 10000.0u 860.347p 0 870.749p 0 870.75p 10000.0u 870.751p 0 882.578p 0 882.579p 10000.0u 882.58p 0 887.993p 0 887.994p 10000.0u 887.995p 0 889.253p 0 889.254p 10000.0u 889.255p 0 910.019p 0 910.02p 10000.0u 910.021p 0 916.697p 0 916.698p 10000.0u 916.699p 0 924.323p 0 924.324p 10000.0u 924.325p 0 932.207p 0 932.208p 10000.0u 932.209p 0 934.322p 0 934.323p 10000.0u 934.324p 0 935.138p 0 935.139p 10000.0u 935.14p 0 965.525p 0 965.526p 10000.0u 965.527p 0 976.724p 0 976.725p 10000.0u 976.726p 0 980.105p 0 980.106p 10000.0u 980.107p 0 985.736p 0 985.737p 10000.0u 985.738p 0 990.632p 0 990.633p 10000.0u 990.634p 0 992.906p 0 992.907p 10000.0u 992.908p 0 995.522p 0 995.523p 10000.0u 995.524p 0)
IIN70 0 71 pwl(0 0 4.619p 0 4.62p 10000.0u 4.621p 0 8.063p 0 8.064p 10000.0u 8.065p 0 8.678p 0 8.679p 10000.0u 8.68p 0 9.362p 0 9.363p 10000.0u 9.364p 0 12.686p 0 12.687p 10000.0u 12.688p 0 32.357p 0 32.358p 10000.0u 32.359p 0 46.274p 0 46.275p 10000.0u 46.276p 0 54.674p 0 54.675p 10000.0u 54.676p 0 59.405p 0 59.406p 10000.0u 59.407p 0 81.974p 0 81.975p 10000.0u 81.976p 0 109.697p 0 109.698p 10000.0u 109.699p 0 118.022p 0 118.023p 10000.0u 118.024p 0 148.163p 0 148.164p 10000.0u 148.165p 0 173.9p 0 173.901p 10000.0u 173.902p 0 179.462p 0 179.463p 10000.0u 179.464p 0 181.577p 0 181.578p 10000.0u 181.579p 0 190.307p 0 190.308p 10000.0u 190.309p 0 193.916p 0 193.917p 10000.0u 193.918p 0 208.142p 0 208.143p 10000.0u 208.144p 0 208.292p 0 208.293p 10000.0u 208.294p 0 216.926p 0 216.927p 10000.0u 216.928p 0 239.441p 0 239.442p 10000.0u 239.443p 0 243.221p 0 243.222p 10000.0u 243.223p 0 247.538p 0 247.539p 10000.0u 247.54p 0 249.818p 0 249.819p 10000.0u 249.82p 0 250.601p 0 250.602p 10000.0u 250.603p 0 251.093p 0 251.094p 10000.0u 251.095p 0 259.772p 0 259.773p 10000.0u 259.774p 0 264.263p 0 264.264p 10000.0u 264.265p 0 272.513p 0 272.514p 10000.0u 272.515p 0 281.861p 0 281.862p 10000.0u 281.863p 0 287.834p 0 287.835p 10000.0u 287.836p 0 294.281p 0 294.282p 10000.0u 294.283p 0 299.924p 0 299.925p 10000.0u 299.926p 0 303.458p 0 303.459p 10000.0u 303.46p 0 330.962p 0 330.963p 10000.0u 330.964p 0 349.622p 0 349.623p 10000.0u 349.624p 0 355.298p 0 355.299p 10000.0u 355.3p 0 371.003p 0 371.004p 10000.0u 371.005p 0 380.888p 0 380.889p 10000.0u 380.89p 0 383.543p 0 383.544p 10000.0u 383.545p 0 391.736p 0 391.737p 10000.0u 391.738p 0 392.882p 0 392.883p 10000.0u 392.884p 0 400.289p 0 400.29p 10000.0u 400.291p 0 414.671p 0 414.672p 10000.0u 414.673p 0 418.745p 0 418.746p 10000.0u 418.747p 0 419.912p 0 419.913p 10000.0u 419.914p 0 425.114p 0 425.115p 10000.0u 425.116p 0 429.161p 0 429.162p 10000.0u 429.163p 0 437.117p 0 437.118p 10000.0u 437.119p 0 442.727p 0 442.728p 10000.0u 442.729p 0 445.889p 0 445.89p 10000.0u 445.891p 0 448.178p 0 448.179p 10000.0u 448.18p 0 449.81p 0 449.811p 10000.0u 449.812p 0 457.01p 0 457.011p 10000.0u 457.012p 0 461.72p 0 461.721p 10000.0u 461.722p 0 467.417p 0 467.418p 10000.0u 467.419p 0 469.058p 0 469.059p 10000.0u 469.06p 0 476.528p 0 476.529p 10000.0u 476.53p 0 476.972p 0 476.973p 10000.0u 476.974p 0 490.076p 0 490.077p 10000.0u 490.078p 0 491.597p 0 491.598p 10000.0u 491.599p 0 500.849p 0 500.85p 10000.0u 500.851p 0 504.926p 0 504.927p 10000.0u 504.928p 0 511.514p 0 511.515p 10000.0u 511.516p 0 513.578p 0 513.579p 10000.0u 513.58p 0 515.06p 0 515.061p 10000.0u 515.062p 0 516.962p 0 516.963p 10000.0u 516.964p 0 517.916p 0 517.917p 10000.0u 517.918p 0 541.577p 0 541.578p 10000.0u 541.579p 0 574.559p 0 574.56p 10000.0u 574.561p 0 577.787p 0 577.788p 10000.0u 577.789p 0 578.612p 0 578.613p 10000.0u 578.614p 0 584.624p 0 584.625p 10000.0u 584.626p 0 589.793p 0 589.794p 10000.0u 589.795p 0 590.075p 0 590.076p 10000.0u 590.077p 0 593.384p 0 593.385p 10000.0u 593.386p 0 600.839p 0 600.84p 10000.0u 600.841p 0 613.085p 0 613.086p 10000.0u 613.087p 0 630.125p 0 630.126p 10000.0u 630.127p 0 648.278p 0 648.279p 10000.0u 648.28p 0 653.564p 0 653.565p 10000.0u 653.566p 0 661.307p 0 661.308p 10000.0u 661.309p 0 683.51p 0 683.511p 10000.0u 683.512p 0 689.648p 0 689.649p 10000.0u 689.65p 0 689.957p 0 689.958p 10000.0u 689.959p 0 690.41p 0 690.411p 10000.0u 690.412p 0 704.447p 0 704.448p 10000.0u 704.449p 0 706.214p 0 706.215p 10000.0u 706.216p 0 730.583p 0 730.584p 10000.0u 730.585p 0 770.084p 0 770.085p 10000.0u 770.086p 0 774.146p 0 774.147p 10000.0u 774.148p 0 783.158p 0 783.159p 10000.0u 783.16p 0 783.965p 0 783.966p 10000.0u 783.967p 0 794.696p 0 794.697p 10000.0u 794.698p 0 802.046p 0 802.047p 10000.0u 802.048p 0 834.746p 0 834.747p 10000.0u 834.748p 0 852.533p 0 852.534p 10000.0u 852.535p 0 854.222p 0 854.223p 10000.0u 854.224p 0 871.445p 0 871.446p 10000.0u 871.447p 0 871.574p 0 871.575p 10000.0u 871.576p 0 879.302p 0 879.303p 10000.0u 879.304p 0 883.952p 0 883.953p 10000.0u 883.954p 0 900.572p 0 900.573p 10000.0u 900.574p 0 910.439p 0 910.44p 10000.0u 910.441p 0 913.247p 0 913.248p 10000.0u 913.249p 0 925.559p 0 925.56p 10000.0u 925.561p 0 926.801p 0 926.802p 10000.0u 926.803p 0 931.328p 0 931.329p 10000.0u 931.33p 0 931.535p 0 931.536p 10000.0u 931.537p 0 939.794p 0 939.795p 10000.0u 939.796p 0 941.786p 0 941.787p 10000.0u 941.788p 0 962.027p 0 962.028p 10000.0u 962.029p 0 977.153p 0 977.154p 10000.0u 977.155p 0 979.916p 0 979.917p 10000.0u 979.918p 0 990.986p 0 990.987p 10000.0u 990.988p 0 999.227p 0 999.228p 10000.0u 999.229p 0)
IIN71 0 72 pwl(0 0 84.26p 0 84.261p 10000.0u 84.262p 0 86.147p 0 86.148p 10000.0u 86.149p 0 86.15p 0 86.151p 10000.0u 86.152p 0 90.29p 0 90.291p 10000.0u 90.292p 0 93.293p 0 93.294p 10000.0u 93.295p 0 133.025p 0 133.026p 10000.0u 133.027p 0 141.542p 0 141.543p 10000.0u 141.544p 0 146.936p 0 146.937p 10000.0u 146.938p 0 152.123p 0 152.124p 10000.0u 152.125p 0 159.332p 0 159.333p 10000.0u 159.334p 0 163.403p 0 163.404p 10000.0u 163.405p 0 172.235p 0 172.236p 10000.0u 172.237p 0 180.743p 0 180.744p 10000.0u 180.745p 0 185.477p 0 185.478p 10000.0u 185.479p 0 187.226p 0 187.227p 10000.0u 187.228p 0 201.554p 0 201.555p 10000.0u 201.556p 0 204.281p 0 204.282p 10000.0u 204.283p 0 211.169p 0 211.17p 10000.0u 211.171p 0 214.352p 0 214.353p 10000.0u 214.354p 0 224.288p 0 224.289p 10000.0u 224.29p 0 244.064p 0 244.065p 10000.0u 244.066p 0 252.383p 0 252.384p 10000.0u 252.385p 0 258.623p 0 258.624p 10000.0u 258.625p 0 285.308p 0 285.309p 10000.0u 285.31p 0 306.479p 0 306.48p 10000.0u 306.481p 0 315.245p 0 315.246p 10000.0u 315.247p 0 328.034p 0 328.035p 10000.0u 328.036p 0 335.342p 0 335.343p 10000.0u 335.344p 0 361.175p 0 361.176p 10000.0u 361.177p 0 388.898p 0 388.899p 10000.0u 388.9p 0 405.68p 0 405.681p 10000.0u 405.682p 0 421.067p 0 421.068p 10000.0u 421.069p 0 426.83p 0 426.831p 10000.0u 426.832p 0 449.651p 0 449.652p 10000.0u 449.653p 0 463.751p 0 463.752p 10000.0u 463.753p 0 482.423p 0 482.424p 10000.0u 482.425p 0 483.605p 0 483.606p 10000.0u 483.607p 0 485.996p 0 485.997p 10000.0u 485.998p 0 495.602p 0 495.603p 10000.0u 495.604p 0 506.327p 0 506.328p 10000.0u 506.329p 0 509.126p 0 509.127p 10000.0u 509.128p 0 513.782p 0 513.783p 10000.0u 513.784p 0 528.656p 0 528.657p 10000.0u 528.658p 0 533.405p 0 533.406p 10000.0u 533.407p 0 549.119p 0 549.12p 10000.0u 549.121p 0 554.372p 0 554.373p 10000.0u 554.374p 0 554.597p 0 554.598p 10000.0u 554.599p 0 572.774p 0 572.775p 10000.0u 572.776p 0 585.035p 0 585.036p 10000.0u 585.037p 0 585.266p 0 585.267p 10000.0u 585.268p 0 589.271p 0 589.272p 10000.0u 589.273p 0 595.355p 0 595.356p 10000.0u 595.357p 0 597.443p 0 597.444p 10000.0u 597.445p 0 598.889p 0 598.89p 10000.0u 598.891p 0 605.654p 0 605.655p 10000.0u 605.656p 0 622.436p 0 622.437p 10000.0u 622.438p 0 636.437p 0 636.438p 10000.0u 636.439p 0 640.136p 0 640.137p 10000.0u 640.138p 0 647.18p 0 647.181p 10000.0u 647.182p 0 648.773p 0 648.774p 10000.0u 648.775p 0 656.753p 0 656.754p 10000.0u 656.755p 0 661.913p 0 661.914p 10000.0u 661.915p 0 662.039p 0 662.04p 10000.0u 662.041p 0 690.128p 0 690.129p 10000.0u 690.13p 0 704.129p 0 704.13p 10000.0u 704.131p 0 731.84p 0 731.841p 10000.0u 731.842p 0 734.222p 0 734.223p 10000.0u 734.224p 0 747.56p 0 747.561p 10000.0u 747.562p 0 752.411p 0 752.412p 10000.0u 752.413p 0 760.601p 0 760.602p 10000.0u 760.603p 0 770.423p 0 770.424p 10000.0u 770.425p 0 771.656p 0 771.657p 10000.0u 771.658p 0 815.774p 0 815.775p 10000.0u 815.776p 0 819.767p 0 819.768p 10000.0u 819.769p 0 831.398p 0 831.399p 10000.0u 831.4p 0 843.395p 0 843.396p 10000.0u 843.397p 0 845.009p 0 845.01p 10000.0u 845.011p 0 848.459p 0 848.46p 10000.0u 848.461p 0 853.673p 0 853.674p 10000.0u 853.675p 0 862.352p 0 862.353p 10000.0u 862.354p 0 863.225p 0 863.226p 10000.0u 863.227p 0 881.255p 0 881.256p 10000.0u 881.257p 0 883.805p 0 883.806p 10000.0u 883.807p 0 889.634p 0 889.635p 10000.0u 889.636p 0 905.315p 0 905.316p 10000.0u 905.317p 0 916.685p 0 916.686p 10000.0u 916.687p 0 924.566p 0 924.567p 10000.0u 924.568p 0 952.559p 0 952.56p 10000.0u 952.561p 0 972.647p 0 972.648p 10000.0u 972.649p 0 973.073p 0 973.074p 10000.0u 973.075p 0 980.261p 0 980.262p 10000.0u 980.263p 0 983.954p 0 983.955p 10000.0u 983.956p 0 985.571p 0 985.572p 10000.0u 985.573p 0 991.907p 0 991.908p 10000.0u 991.909p 0)
IIN72 0 73 pwl(0 0 1.853p 0 1.854p 10000.0u 1.855p 0 6.389p 0 6.39p 10000.0u 6.391p 0 13.337p 0 13.338p 10000.0u 13.339p 0 13.931p 0 13.932p 10000.0u 13.933p 0 18.302p 0 18.303p 10000.0u 18.304p 0 25.355p 0 25.356p 10000.0u 25.357p 0 25.817p 0 25.818p 10000.0u 25.819p 0 27.323p 0 27.324p 10000.0u 27.325p 0 44.774p 0 44.775p 10000.0u 44.776p 0 53.159p 0 53.16p 10000.0u 53.161p 0 54.512p 0 54.513p 10000.0u 54.514p 0 63.704p 0 63.705p 10000.0u 63.706p 0 63.764p 0 63.765p 10000.0u 63.766p 0 71.099p 0 71.1p 10000.0u 71.101p 0 101.087p 0 101.088p 10000.0u 101.089p 0 112.022p 0 112.023p 10000.0u 112.024p 0 120.872p 0 120.873p 10000.0u 120.874p 0 121.7p 0 121.701p 10000.0u 121.702p 0 124.355p 0 124.356p 10000.0u 124.357p 0 127.94p 0 127.941p 10000.0u 127.942p 0 138.698p 0 138.699p 10000.0u 138.7p 0 151.826p 0 151.827p 10000.0u 151.828p 0 154.007p 0 154.008p 10000.0u 154.009p 0 172.214p 0 172.215p 10000.0u 172.216p 0 188.285p 0 188.286p 10000.0u 188.287p 0 188.666p 0 188.667p 10000.0u 188.668p 0 195.098p 0 195.099p 10000.0u 195.1p 0 207.341p 0 207.342p 10000.0u 207.343p 0 216.014p 0 216.015p 10000.0u 216.016p 0 225.974p 0 225.975p 10000.0u 225.976p 0 235.571p 0 235.572p 10000.0u 235.573p 0 235.952p 0 235.953p 10000.0u 235.954p 0 242.174p 0 242.175p 10000.0u 242.176p 0 269.744p 0 269.745p 10000.0u 269.746p 0 271.46p 0 271.461p 10000.0u 271.462p 0 289.529p 0 289.53p 10000.0u 289.531p 0 313.52p 0 313.521p 10000.0u 313.522p 0 333.128p 0 333.129p 10000.0u 333.13p 0 335.594p 0 335.595p 10000.0u 335.596p 0 349.946p 0 349.947p 10000.0u 349.948p 0 350.414p 0 350.415p 10000.0u 350.416p 0 356.744p 0 356.745p 10000.0u 356.746p 0 368.903p 0 368.904p 10000.0u 368.905p 0 384.272p 0 384.273p 10000.0u 384.274p 0 388.967p 0 388.968p 10000.0u 388.969p 0 391.694p 0 391.695p 10000.0u 391.696p 0 395.822p 0 395.823p 10000.0u 395.824p 0 405.008p 0 405.009p 10000.0u 405.01p 0 409.595p 0 409.596p 10000.0u 409.597p 0 447.539p 0 447.54p 10000.0u 447.541p 0 465.53p 0 465.531p 10000.0u 465.532p 0 466.304p 0 466.305p 10000.0u 466.306p 0 484.475p 0 484.476p 10000.0u 484.477p 0 499.649p 0 499.65p 10000.0u 499.651p 0 518.66p 0 518.661p 10000.0u 518.662p 0 525.764p 0 525.765p 10000.0u 525.766p 0 533.048p 0 533.049p 10000.0u 533.05p 0 558.593p 0 558.594p 10000.0u 558.595p 0 566.555p 0 566.556p 10000.0u 566.557p 0 572.933p 0 572.934p 10000.0u 572.935p 0 580.943p 0 580.944p 10000.0u 580.945p 0 591.116p 0 591.117p 10000.0u 591.118p 0 598.31p 0 598.311p 10000.0u 598.312p 0 600.695p 0 600.696p 10000.0u 600.697p 0 620.873p 0 620.874p 10000.0u 620.875p 0 633.2p 0 633.201p 10000.0u 633.202p 0 634.595p 0 634.596p 10000.0u 634.597p 0 650.174p 0 650.175p 10000.0u 650.176p 0 659.426p 0 659.427p 10000.0u 659.428p 0 681.227p 0 681.228p 10000.0u 681.229p 0 682.103p 0 682.104p 10000.0u 682.105p 0 708.203p 0 708.204p 10000.0u 708.205p 0 715.484p 0 715.485p 10000.0u 715.486p 0 716.606p 0 716.607p 10000.0u 716.608p 0 741.872p 0 741.873p 10000.0u 741.874p 0 748.448p 0 748.449p 10000.0u 748.45p 0 750.143p 0 750.144p 10000.0u 750.145p 0 775.973p 0 775.974p 10000.0u 775.975p 0 778.07p 0 778.071p 10000.0u 778.072p 0 814.919p 0 814.92p 10000.0u 814.921p 0 821.501p 0 821.502p 10000.0u 821.503p 0 838.979p 0 838.98p 10000.0u 838.981p 0 852.962p 0 852.963p 10000.0u 852.964p 0 863.975p 0 863.976p 10000.0u 863.977p 0 866.912p 0 866.913p 10000.0u 866.914p 0 890.099p 0 890.1p 10000.0u 890.101p 0 891.095p 0 891.096p 10000.0u 891.097p 0 895.04p 0 895.041p 10000.0u 895.042p 0 907.649p 0 907.65p 10000.0u 907.651p 0 908.909p 0 908.91p 10000.0u 908.911p 0 912.446p 0 912.447p 10000.0u 912.448p 0 932.261p 0 932.262p 10000.0u 932.263p 0 932.945p 0 932.946p 10000.0u 932.947p 0 933.281p 0 933.282p 10000.0u 933.283p 0 938.438p 0 938.439p 10000.0u 938.44p 0 940.955p 0 940.956p 10000.0u 940.957p 0 942.275p 0 942.276p 10000.0u 942.277p 0 956.144p 0 956.145p 10000.0u 956.146p 0 964.568p 0 964.569p 10000.0u 964.57p 0 969.116p 0 969.117p 10000.0u 969.118p 0)
IIN73 0 74 pwl(0 0 3.446p 0 3.447p 10000.0u 3.448p 0 7.034p 0 7.035p 10000.0u 7.036p 0 10.667p 0 10.668p 10000.0u 10.669p 0 15.119p 0 15.12p 10000.0u 15.121p 0 27.125p 0 27.126p 10000.0u 27.127p 0 41.774p 0 41.775p 10000.0u 41.776p 0 54.674p 0 54.675p 10000.0u 54.676p 0 64.772p 0 64.773p 10000.0u 64.774p 0 84.425p 0 84.426p 10000.0u 84.427p 0 85.25p 0 85.251p 10000.0u 85.252p 0 95.093p 0 95.094p 10000.0u 95.095p 0 103.454p 0 103.455p 10000.0u 103.456p 0 107.975p 0 107.976p 10000.0u 107.977p 0 108.236p 0 108.237p 10000.0u 108.238p 0 131.12p 0 131.121p 10000.0u 131.122p 0 137.945p 0 137.946p 10000.0u 137.947p 0 141.767p 0 141.768p 10000.0u 141.769p 0 153.362p 0 153.363p 10000.0u 153.364p 0 168.578p 0 168.579p 10000.0u 168.58p 0 175.856p 0 175.857p 10000.0u 175.858p 0 177.545p 0 177.546p 10000.0u 177.547p 0 187.04p 0 187.041p 10000.0u 187.042p 0 189.626p 0 189.627p 10000.0u 189.628p 0 204.239p 0 204.24p 10000.0u 204.241p 0 223.814p 0 223.815p 10000.0u 223.816p 0 239.873p 0 239.874p 10000.0u 239.875p 0 239.972p 0 239.973p 10000.0u 239.974p 0 251.045p 0 251.046p 10000.0u 251.047p 0 252.755p 0 252.756p 10000.0u 252.757p 0 260.462p 0 260.463p 10000.0u 260.464p 0 279.308p 0 279.309p 10000.0u 279.31p 0 301.388p 0 301.389p 10000.0u 301.39p 0 330.5p 0 330.501p 10000.0u 330.502p 0 336.752p 0 336.753p 10000.0u 336.754p 0 344.069p 0 344.07p 10000.0u 344.071p 0 356.024p 0 356.025p 10000.0u 356.026p 0 361.136p 0 361.137p 10000.0u 361.138p 0 362.681p 0 362.682p 10000.0u 362.683p 0 387.626p 0 387.627p 10000.0u 387.628p 0 389.837p 0 389.838p 10000.0u 389.839p 0 401.726p 0 401.727p 10000.0u 401.728p 0 408.116p 0 408.117p 10000.0u 408.118p 0 417.833p 0 417.834p 10000.0u 417.835p 0 429.653p 0 429.654p 10000.0u 429.655p 0 430.655p 0 430.656p 10000.0u 430.657p 0 432.377p 0 432.378p 10000.0u 432.379p 0 459.44p 0 459.441p 10000.0u 459.442p 0 474.92p 0 474.921p 10000.0u 474.922p 0 478.001p 0 478.002p 10000.0u 478.003p 0 494.63p 0 494.631p 10000.0u 494.632p 0 494.651p 0 494.652p 10000.0u 494.653p 0 500.402p 0 500.403p 10000.0u 500.404p 0 505.427p 0 505.428p 10000.0u 505.429p 0 535.613p 0 535.614p 10000.0u 535.615p 0 537.824p 0 537.825p 10000.0u 537.826p 0 542.63p 0 542.631p 10000.0u 542.632p 0 563.177p 0 563.178p 10000.0u 563.179p 0 568.091p 0 568.092p 10000.0u 568.093p 0 578.804p 0 578.805p 10000.0u 578.806p 0 589.238p 0 589.239p 10000.0u 589.24p 0 592.91p 0 592.911p 10000.0u 592.912p 0 593.906p 0 593.907p 10000.0u 593.908p 0 598.004p 0 598.005p 10000.0u 598.006p 0 614.03p 0 614.031p 10000.0u 614.032p 0 617.522p 0 617.523p 10000.0u 617.524p 0 621.962p 0 621.963p 10000.0u 621.964p 0 632.414p 0 632.415p 10000.0u 632.416p 0 634.013p 0 634.014p 10000.0u 634.015p 0 642.65p 0 642.651p 10000.0u 642.652p 0 643.937p 0 643.938p 10000.0u 643.939p 0 678.026p 0 678.027p 10000.0u 678.028p 0 704.354p 0 704.355p 10000.0u 704.356p 0 707.459p 0 707.46p 10000.0u 707.461p 0 712.928p 0 712.929p 10000.0u 712.93p 0 721.013p 0 721.014p 10000.0u 721.015p 0 726.029p 0 726.03p 10000.0u 726.031p 0 732.869p 0 732.87p 10000.0u 732.871p 0 738.329p 0 738.33p 10000.0u 738.331p 0 770.621p 0 770.622p 10000.0u 770.623p 0 772.508p 0 772.509p 10000.0u 772.51p 0 773.372p 0 773.373p 10000.0u 773.374p 0 786.908p 0 786.909p 10000.0u 786.91p 0 792.149p 0 792.15p 10000.0u 792.151p 0 793.676p 0 793.677p 10000.0u 793.678p 0 794.171p 0 794.172p 10000.0u 794.173p 0 806.666p 0 806.667p 10000.0u 806.668p 0 843.134p 0 843.135p 10000.0u 843.136p 0 857.852p 0 857.853p 10000.0u 857.854p 0 862.529p 0 862.53p 10000.0u 862.531p 0 896.729p 0 896.73p 10000.0u 896.731p 0 897.95p 0 897.951p 10000.0u 897.952p 0 903.737p 0 903.738p 10000.0u 903.739p 0 913.292p 0 913.293p 10000.0u 913.294p 0 921.071p 0 921.072p 10000.0u 921.073p 0 922.559p 0 922.56p 10000.0u 922.561p 0 925.907p 0 925.908p 10000.0u 925.909p 0 928.82p 0 928.821p 10000.0u 928.822p 0 933.209p 0 933.21p 10000.0u 933.211p 0 946.319p 0 946.32p 10000.0u 946.321p 0 949.961p 0 949.962p 10000.0u 949.963p 0 950.435p 0 950.436p 10000.0u 950.437p 0 951.767p 0 951.768p 10000.0u 951.769p 0 952.283p 0 952.284p 10000.0u 952.285p 0 978.956p 0 978.957p 10000.0u 978.958p 0 981.122p 0 981.123p 10000.0u 981.124p 0 988.412p 0 988.413p 10000.0u 988.414p 0 994.607p 0 994.608p 10000.0u 994.609p 0)
IIN74 0 75 pwl(0 0 15.209p 0 15.21p 10000.0u 15.211p 0 26.639p 0 26.64p 10000.0u 26.641p 0 42.245p 0 42.246p 10000.0u 42.247p 0 43.13p 0 43.131p 10000.0u 43.132p 0 47.249p 0 47.25p 10000.0u 47.251p 0 63.122p 0 63.123p 10000.0u 63.124p 0 77.153p 0 77.154p 10000.0u 77.155p 0 86.177p 0 86.178p 10000.0u 86.179p 0 87.353p 0 87.354p 10000.0u 87.355p 0 100.892p 0 100.893p 10000.0u 100.894p 0 100.994p 0 100.995p 10000.0u 100.996p 0 124.076p 0 124.077p 10000.0u 124.078p 0 136.448p 0 136.449p 10000.0u 136.45p 0 166.106p 0 166.107p 10000.0u 166.108p 0 178.616p 0 178.617p 10000.0u 178.618p 0 185.438p 0 185.439p 10000.0u 185.44p 0 233.372p 0 233.373p 10000.0u 233.374p 0 235.211p 0 235.212p 10000.0u 235.213p 0 250.412p 0 250.413p 10000.0u 250.414p 0 252.977p 0 252.978p 10000.0u 252.979p 0 258.896p 0 258.897p 10000.0u 258.898p 0 278.678p 0 278.679p 10000.0u 278.68p 0 291.719p 0 291.72p 10000.0u 291.721p 0 302.957p 0 302.958p 10000.0u 302.959p 0 324.182p 0 324.183p 10000.0u 324.184p 0 332.396p 0 332.397p 10000.0u 332.398p 0 336.548p 0 336.549p 10000.0u 336.55p 0 355.829p 0 355.83p 10000.0u 355.831p 0 369.545p 0 369.546p 10000.0u 369.547p 0 372.158p 0 372.159p 10000.0u 372.16p 0 380.165p 0 380.166p 10000.0u 380.167p 0 381.074p 0 381.075p 10000.0u 381.076p 0 409.637p 0 409.638p 10000.0u 409.639p 0 410.021p 0 410.022p 10000.0u 410.023p 0 411.419p 0 411.42p 10000.0u 411.421p 0 411.533p 0 411.534p 10000.0u 411.535p 0 444.941p 0 444.942p 10000.0u 444.943p 0 453.398p 0 453.399p 10000.0u 453.4p 0 465.128p 0 465.129p 10000.0u 465.13p 0 492.698p 0 492.699p 10000.0u 492.7p 0 503.768p 0 503.769p 10000.0u 503.77p 0 514.007p 0 514.008p 10000.0u 514.009p 0 515.447p 0 515.448p 10000.0u 515.449p 0 518.213p 0 518.214p 10000.0u 518.215p 0 542.042p 0 542.043p 10000.0u 542.044p 0 557.546p 0 557.547p 10000.0u 557.548p 0 570.542p 0 570.543p 10000.0u 570.544p 0 600.968p 0 600.969p 10000.0u 600.97p 0 603.008p 0 603.009p 10000.0u 603.01p 0 609.98p 0 609.981p 10000.0u 609.982p 0 610.496p 0 610.497p 10000.0u 610.498p 0 621.989p 0 621.99p 10000.0u 621.991p 0 626.216p 0 626.217p 10000.0u 626.218p 0 628.955p 0 628.956p 10000.0u 628.957p 0 629.303p 0 629.304p 10000.0u 629.305p 0 642.506p 0 642.507p 10000.0u 642.508p 0 673.937p 0 673.938p 10000.0u 673.939p 0 679.286p 0 679.287p 10000.0u 679.288p 0 691.676p 0 691.677p 10000.0u 691.678p 0 699.065p 0 699.066p 10000.0u 699.067p 0 714.962p 0 714.963p 10000.0u 714.964p 0 720.395p 0 720.396p 10000.0u 720.397p 0 746.489p 0 746.49p 10000.0u 746.491p 0 756.191p 0 756.192p 10000.0u 756.193p 0 759.905p 0 759.906p 10000.0u 759.907p 0 790.667p 0 790.668p 10000.0u 790.669p 0 793.433p 0 793.434p 10000.0u 793.435p 0 796.145p 0 796.146p 10000.0u 796.147p 0 815.057p 0 815.058p 10000.0u 815.059p 0 819.485p 0 819.486p 10000.0u 819.487p 0 828.773p 0 828.774p 10000.0u 828.775p 0 846.023p 0 846.024p 10000.0u 846.025p 0 851.273p 0 851.274p 10000.0u 851.275p 0 860.507p 0 860.508p 10000.0u 860.509p 0 861.965p 0 861.966p 10000.0u 861.967p 0 862.604p 0 862.605p 10000.0u 862.606p 0 878.909p 0 878.91p 10000.0u 878.911p 0 891.281p 0 891.282p 10000.0u 891.283p 0 891.791p 0 891.792p 10000.0u 891.793p 0 895.745p 0 895.746p 10000.0u 895.747p 0 911.894p 0 911.895p 10000.0u 911.896p 0 913.43p 0 913.431p 10000.0u 913.432p 0 929.123p 0 929.124p 10000.0u 929.125p 0 929.48p 0 929.481p 10000.0u 929.482p 0 963.713p 0 963.714p 10000.0u 963.715p 0 964.574p 0 964.575p 10000.0u 964.576p 0 966.194p 0 966.195p 10000.0u 966.196p 0)
IIN75 0 76 pwl(0 0 7.337p 0 7.338p 10000.0u 7.339p 0 26.378p 0 26.379p 10000.0u 26.38p 0 38.033p 0 38.034p 10000.0u 38.035p 0 40.274p 0 40.275p 10000.0u 40.276p 0 65.762p 0 65.763p 10000.0u 65.764p 0 72.176p 0 72.177p 10000.0u 72.178p 0 73.652p 0 73.653p 10000.0u 73.654p 0 74.807p 0 74.808p 10000.0u 74.809p 0 78.542p 0 78.543p 10000.0u 78.544p 0 102.224p 0 102.225p 10000.0u 102.226p 0 105.659p 0 105.66p 10000.0u 105.661p 0 106.07p 0 106.071p 10000.0u 106.072p 0 131.042p 0 131.043p 10000.0u 131.044p 0 148.334p 0 148.335p 10000.0u 148.336p 0 148.478p 0 148.479p 10000.0u 148.48p 0 156.59p 0 156.591p 10000.0u 156.592p 0 162.26p 0 162.261p 10000.0u 162.262p 0 164.924p 0 164.925p 10000.0u 164.926p 0 218.387p 0 218.388p 10000.0u 218.389p 0 222.182p 0 222.183p 10000.0u 222.184p 0 224.327p 0 224.328p 10000.0u 224.329p 0 234.305p 0 234.306p 10000.0u 234.307p 0 252.548p 0 252.549p 10000.0u 252.55p 0 261.464p 0 261.465p 10000.0u 261.466p 0 286.253p 0 286.254p 10000.0u 286.255p 0 320.285p 0 320.286p 10000.0u 320.287p 0 370.418p 0 370.419p 10000.0u 370.42p 0 378.863p 0 378.864p 10000.0u 378.865p 0 380.099p 0 380.1p 10000.0u 380.101p 0 392.708p 0 392.709p 10000.0u 392.71p 0 412.31p 0 412.311p 10000.0u 412.312p 0 416.255p 0 416.256p 10000.0u 416.257p 0 417.419p 0 417.42p 10000.0u 417.421p 0 428.855p 0 428.856p 10000.0u 428.857p 0 433.427p 0 433.428p 10000.0u 433.429p 0 436.061p 0 436.062p 10000.0u 436.063p 0 436.73p 0 436.731p 10000.0u 436.732p 0 447.755p 0 447.756p 10000.0u 447.757p 0 458.465p 0 458.466p 10000.0u 458.467p 0 460.049p 0 460.05p 10000.0u 460.051p 0 465.911p 0 465.912p 10000.0u 465.913p 0 468.938p 0 468.939p 10000.0u 468.94p 0 472.805p 0 472.806p 10000.0u 472.807p 0 487.058p 0 487.059p 10000.0u 487.06p 0 497.525p 0 497.526p 10000.0u 497.527p 0 508.193p 0 508.194p 10000.0u 508.195p 0 510.581p 0 510.582p 10000.0u 510.583p 0 513.923p 0 513.924p 10000.0u 513.925p 0 535.841p 0 535.842p 10000.0u 535.843p 0 538.202p 0 538.203p 10000.0u 538.204p 0 538.517p 0 538.518p 10000.0u 538.519p 0 552.086p 0 552.087p 10000.0u 552.088p 0 556.265p 0 556.266p 10000.0u 556.267p 0 568.094p 0 568.095p 10000.0u 568.096p 0 574.496p 0 574.497p 10000.0u 574.498p 0 578.903p 0 578.904p 10000.0u 578.905p 0 598.139p 0 598.14p 10000.0u 598.141p 0 610.235p 0 610.236p 10000.0u 610.237p 0 610.958p 0 610.959p 10000.0u 610.96p 0 620.75p 0 620.751p 10000.0u 620.752p 0 622.094p 0 622.095p 10000.0u 622.096p 0 636.731p 0 636.732p 10000.0u 636.733p 0 644.534p 0 644.535p 10000.0u 644.536p 0 656.972p 0 656.973p 10000.0u 656.974p 0 665.831p 0 665.832p 10000.0u 665.833p 0 667.805p 0 667.806p 10000.0u 667.807p 0 668.237p 0 668.238p 10000.0u 668.239p 0 677.987p 0 677.988p 10000.0u 677.989p 0 689.603p 0 689.604p 10000.0u 689.605p 0 695.651p 0 695.652p 10000.0u 695.653p 0 716.774p 0 716.775p 10000.0u 716.776p 0 725.357p 0 725.358p 10000.0u 725.359p 0 730.829p 0 730.83p 10000.0u 730.831p 0 747.806p 0 747.807p 10000.0u 747.808p 0 752.087p 0 752.088p 10000.0u 752.089p 0 761.249p 0 761.25p 10000.0u 761.251p 0 764.747p 0 764.748p 10000.0u 764.749p 0 769.949p 0 769.95p 10000.0u 769.951p 0 785.558p 0 785.559p 10000.0u 785.56p 0 794.72p 0 794.721p 10000.0u 794.722p 0 794.954p 0 794.955p 10000.0u 794.956p 0 812.516p 0 812.517p 10000.0u 812.518p 0 817.886p 0 817.887p 10000.0u 817.888p 0 829.769p 0 829.77p 10000.0u 829.771p 0 855.137p 0 855.138p 10000.0u 855.139p 0 864.656p 0 864.657p 10000.0u 864.658p 0 865.607p 0 865.608p 10000.0u 865.609p 0 874.889p 0 874.89p 10000.0u 874.891p 0 888.338p 0 888.339p 10000.0u 888.34p 0 890.231p 0 890.232p 10000.0u 890.233p 0 892.277p 0 892.278p 10000.0u 892.279p 0 897.185p 0 897.186p 10000.0u 897.187p 0 901.58p 0 901.581p 10000.0u 901.582p 0 905.177p 0 905.178p 10000.0u 905.179p 0 912.584p 0 912.585p 10000.0u 912.586p 0 912.878p 0 912.879p 10000.0u 912.88p 0 927.437p 0 927.438p 10000.0u 927.439p 0 930.239p 0 930.24p 10000.0u 930.241p 0 930.974p 0 930.975p 10000.0u 930.976p 0 931.934p 0 931.935p 10000.0u 931.936p 0 935.816p 0 935.817p 10000.0u 935.818p 0 939.839p 0 939.84p 10000.0u 939.841p 0 947.03p 0 947.031p 10000.0u 947.032p 0 951.044p 0 951.045p 10000.0u 951.046p 0 995.201p 0 995.202p 10000.0u 995.203p 0)
IIN76 0 77 pwl(0 0 6.743p 0 6.744p 10000.0u 6.745p 0 23.957p 0 23.958p 10000.0u 23.959p 0 24.389p 0 24.39p 10000.0u 24.391p 0 27.266p 0 27.267p 10000.0u 27.268p 0 107.342p 0 107.343p 10000.0u 107.344p 0 112.148p 0 112.149p 10000.0u 112.15p 0 112.892p 0 112.893p 10000.0u 112.894p 0 113.129p 0 113.13p 10000.0u 113.131p 0 135.734p 0 135.735p 10000.0u 135.736p 0 136.844p 0 136.845p 10000.0u 136.846p 0 137.957p 0 137.958p 10000.0u 137.959p 0 175.217p 0 175.218p 10000.0u 175.219p 0 178.388p 0 178.389p 10000.0u 178.39p 0 179.585p 0 179.586p 10000.0u 179.587p 0 199.331p 0 199.332p 10000.0u 199.333p 0 212.882p 0 212.883p 10000.0u 212.884p 0 219.248p 0 219.249p 10000.0u 219.25p 0 230.228p 0 230.229p 10000.0u 230.23p 0 242.252p 0 242.253p 10000.0u 242.254p 0 244.289p 0 244.29p 10000.0u 244.291p 0 253.286p 0 253.287p 10000.0u 253.288p 0 259.268p 0 259.269p 10000.0u 259.27p 0 293.351p 0 293.352p 10000.0u 293.353p 0 303.998p 0 303.999p 10000.0u 304.0p 0 309.506p 0 309.507p 10000.0u 309.508p 0 314.24p 0 314.241p 10000.0u 314.242p 0 318.875p 0 318.876p 10000.0u 318.877p 0 334.886p 0 334.887p 10000.0u 334.888p 0 340.46p 0 340.461p 10000.0u 340.462p 0 344.66p 0 344.661p 10000.0u 344.662p 0 353.276p 0 353.277p 10000.0u 353.278p 0 355.013p 0 355.014p 10000.0u 355.015p 0 362.174p 0 362.175p 10000.0u 362.176p 0 367.067p 0 367.068p 10000.0u 367.069p 0 378.854p 0 378.855p 10000.0u 378.856p 0 388.046p 0 388.047p 10000.0u 388.048p 0 392.231p 0 392.232p 10000.0u 392.233p 0 401.933p 0 401.934p 10000.0u 401.935p 0 404.597p 0 404.598p 10000.0u 404.599p 0 409.442p 0 409.443p 10000.0u 409.444p 0 439.427p 0 439.428p 10000.0u 439.429p 0 439.895p 0 439.896p 10000.0u 439.897p 0 445.784p 0 445.785p 10000.0u 445.786p 0 471.956p 0 471.957p 10000.0u 471.958p 0 478.799p 0 478.8p 10000.0u 478.801p 0 483.908p 0 483.909p 10000.0u 483.91p 0 484.058p 0 484.059p 10000.0u 484.06p 0 486.296p 0 486.297p 10000.0u 486.298p 0 491.84p 0 491.841p 10000.0u 491.842p 0 500.975p 0 500.976p 10000.0u 500.977p 0 523.088p 0 523.089p 10000.0u 523.09p 0 532.208p 0 532.209p 10000.0u 532.21p 0 558.875p 0 558.876p 10000.0u 558.877p 0 565.07p 0 565.071p 10000.0u 565.072p 0 565.244p 0 565.245p 10000.0u 565.246p 0 572.192p 0 572.193p 10000.0u 572.194p 0 572.27p 0 572.271p 10000.0u 572.272p 0 579.941p 0 579.942p 10000.0u 579.943p 0 583.118p 0 583.119p 10000.0u 583.12p 0 601.586p 0 601.587p 10000.0u 601.588p 0 604.004p 0 604.005p 10000.0u 604.006p 0 646.961p 0 646.962p 10000.0u 646.963p 0 648.665p 0 648.666p 10000.0u 648.667p 0 655.091p 0 655.092p 10000.0u 655.093p 0 681.878p 0 681.879p 10000.0u 681.88p 0 694.736p 0 694.737p 10000.0u 694.738p 0 704.444p 0 704.445p 10000.0u 704.446p 0 706.439p 0 706.44p 10000.0u 706.441p 0 729.476p 0 729.477p 10000.0u 729.478p 0 731.417p 0 731.418p 10000.0u 731.419p 0 731.885p 0 731.886p 10000.0u 731.887p 0 741.443p 0 741.444p 10000.0u 741.445p 0 743.285p 0 743.286p 10000.0u 743.287p 0 750.878p 0 750.879p 10000.0u 750.88p 0 781.667p 0 781.668p 10000.0u 781.669p 0 784.253p 0 784.254p 10000.0u 784.255p 0 784.673p 0 784.674p 10000.0u 784.675p 0 787.178p 0 787.179p 10000.0u 787.18p 0 793.697p 0 793.698p 10000.0u 793.699p 0 803.111p 0 803.112p 10000.0u 803.113p 0 806.525p 0 806.526p 10000.0u 806.527p 0 810.341p 0 810.342p 10000.0u 810.343p 0 837.146p 0 837.147p 10000.0u 837.148p 0 861.545p 0 861.546p 10000.0u 861.547p 0 864.035p 0 864.036p 10000.0u 864.037p 0 890.636p 0 890.637p 10000.0u 890.638p 0 891.197p 0 891.198p 10000.0u 891.199p 0 902.135p 0 902.136p 10000.0u 902.137p 0 906.797p 0 906.798p 10000.0u 906.799p 0 928.367p 0 928.368p 10000.0u 928.369p 0 929.426p 0 929.427p 10000.0u 929.428p 0 931.118p 0 931.119p 10000.0u 931.12p 0 956.657p 0 956.658p 10000.0u 956.659p 0 959.627p 0 959.628p 10000.0u 959.629p 0 966.269p 0 966.27p 10000.0u 966.271p 0 966.875p 0 966.876p 10000.0u 966.877p 0 976.751p 0 976.752p 10000.0u 976.753p 0 979.265p 0 979.266p 10000.0u 979.267p 0 986.24p 0 986.241p 10000.0u 986.242p 0 998.996p 0 998.997p 10000.0u 998.998p 0)
IIN77 0 78 pwl(0 0 13.331p 0 13.332p 10000.0u 13.333p 0 14.282p 0 14.283p 10000.0u 14.284p 0 24.914p 0 24.915p 10000.0u 24.916p 0 29.66p 0 29.661p 10000.0u 29.662p 0 33.422p 0 33.423p 10000.0u 33.424p 0 61.1p 0 61.101p 10000.0u 61.102p 0 71.198p 0 71.199p 10000.0u 71.2p 0 99.677p 0 99.678p 10000.0u 99.679p 0 120.146p 0 120.147p 10000.0u 120.148p 0 133.361p 0 133.362p 10000.0u 133.363p 0 142.904p 0 142.905p 10000.0u 142.906p 0 197.543p 0 197.544p 10000.0u 197.545p 0 201.308p 0 201.309p 10000.0u 201.31p 0 209.063p 0 209.064p 10000.0u 209.065p 0 237.575p 0 237.576p 10000.0u 237.577p 0 239.651p 0 239.652p 10000.0u 239.653p 0 239.69p 0 239.691p 10000.0u 239.692p 0 252.314p 0 252.315p 10000.0u 252.316p 0 253.337p 0 253.338p 10000.0u 253.339p 0 261.32p 0 261.321p 10000.0u 261.322p 0 266.528p 0 266.529p 10000.0u 266.53p 0 276.83p 0 276.831p 10000.0u 276.832p 0 279.788p 0 279.789p 10000.0u 279.79p 0 280.49p 0 280.491p 10000.0u 280.492p 0 280.994p 0 280.995p 10000.0u 280.996p 0 281.528p 0 281.529p 10000.0u 281.53p 0 288.47p 0 288.471p 10000.0u 288.472p 0 300.788p 0 300.789p 10000.0u 300.79p 0 312.197p 0 312.198p 10000.0u 312.199p 0 323.735p 0 323.736p 10000.0u 323.737p 0 326.051p 0 326.052p 10000.0u 326.053p 0 340.913p 0 340.914p 10000.0u 340.915p 0 357.443p 0 357.444p 10000.0u 357.445p 0 366.551p 0 366.552p 10000.0u 366.553p 0 373.421p 0 373.422p 10000.0u 373.423p 0 403.886p 0 403.887p 10000.0u 403.888p 0 413.609p 0 413.61p 10000.0u 413.611p 0 425.942p 0 425.943p 10000.0u 425.944p 0 429.728p 0 429.729p 10000.0u 429.73p 0 439.55p 0 439.551p 10000.0u 439.552p 0 443.303p 0 443.304p 10000.0u 443.305p 0 449.225p 0 449.226p 10000.0u 449.227p 0 451.613p 0 451.614p 10000.0u 451.615p 0 452.636p 0 452.637p 10000.0u 452.638p 0 452.693p 0 452.694p 10000.0u 452.695p 0 458.921p 0 458.922p 10000.0u 458.923p 0 470.162p 0 470.163p 10000.0u 470.164p 0 472.43p 0 472.431p 10000.0u 472.432p 0 491.426p 0 491.427p 10000.0u 491.428p 0 519.872p 0 519.873p 10000.0u 519.874p 0 536.72p 0 536.721p 10000.0u 536.722p 0 549.008p 0 549.009p 10000.0u 549.01p 0 557.813p 0 557.814p 10000.0u 557.815p 0 570.218p 0 570.219p 10000.0u 570.22p 0 570.887p 0 570.888p 10000.0u 570.889p 0 573.566p 0 573.567p 10000.0u 573.568p 0 579.092p 0 579.093p 10000.0u 579.094p 0 613.121p 0 613.122p 10000.0u 613.123p 0 625.721p 0 625.722p 10000.0u 625.723p 0 634.724p 0 634.725p 10000.0u 634.726p 0 648.494p 0 648.495p 10000.0u 648.496p 0 662.861p 0 662.862p 10000.0u 662.863p 0 667.22p 0 667.221p 10000.0u 667.222p 0 675.779p 0 675.78p 10000.0u 675.781p 0 676.685p 0 676.686p 10000.0u 676.687p 0 678.269p 0 678.27p 10000.0u 678.271p 0 706.856p 0 706.857p 10000.0u 706.858p 0 716.9p 0 716.901p 10000.0u 716.902p 0 722.063p 0 722.064p 10000.0u 722.065p 0 741.227p 0 741.228p 10000.0u 741.229p 0 746.807p 0 746.808p 10000.0u 746.809p 0 750.641p 0 750.642p 10000.0u 750.643p 0 772.838p 0 772.839p 10000.0u 772.84p 0 785.657p 0 785.658p 10000.0u 785.659p 0 794.468p 0 794.469p 10000.0u 794.47p 0 804.38p 0 804.381p 10000.0u 804.382p 0 818.828p 0 818.829p 10000.0u 818.83p 0 828.857p 0 828.858p 10000.0u 828.859p 0 831.038p 0 831.039p 10000.0u 831.04p 0 833.345p 0 833.346p 10000.0u 833.347p 0 857.588p 0 857.589p 10000.0u 857.59p 0 862.238p 0 862.239p 10000.0u 862.24p 0 887.693p 0 887.694p 10000.0u 887.695p 0 889.964p 0 889.965p 10000.0u 889.966p 0 896.516p 0 896.517p 10000.0u 896.518p 0 908.009p 0 908.01p 10000.0u 908.011p 0 911.993p 0 911.994p 10000.0u 911.995p 0 920.417p 0 920.418p 10000.0u 920.419p 0 929.864p 0 929.865p 10000.0u 929.866p 0 956.168p 0 956.169p 10000.0u 956.17p 0 966.158p 0 966.159p 10000.0u 966.16p 0 974.138p 0 974.139p 10000.0u 974.14p 0 980.507p 0 980.508p 10000.0u 980.509p 0 995.744p 0 995.745p 10000.0u 995.746p 0)
IIN78 0 79 pwl(0 0 38.267p 0 38.268p 10000.0u 38.269p 0 52.115p 0 52.116p 10000.0u 52.117p 0 59.315p 0 59.316p 10000.0u 59.317p 0 76.043p 0 76.044p 10000.0u 76.045p 0 76.157p 0 76.158p 10000.0u 76.159p 0 88.727p 0 88.728p 10000.0u 88.729p 0 96.002p 0 96.003p 10000.0u 96.004p 0 103.562p 0 103.563p 10000.0u 103.564p 0 108.482p 0 108.483p 10000.0u 108.484p 0 136.769p 0 136.77p 10000.0u 136.771p 0 148.409p 0 148.41p 10000.0u 148.411p 0 149.273p 0 149.274p 10000.0u 149.275p 0 149.6p 0 149.601p 10000.0u 149.602p 0 151.703p 0 151.704p 10000.0u 151.705p 0 179.285p 0 179.286p 10000.0u 179.287p 0 195.404p 0 195.405p 10000.0u 195.406p 0 196.01p 0 196.011p 10000.0u 196.012p 0 209.321p 0 209.322p 10000.0u 209.323p 0 211.106p 0 211.107p 10000.0u 211.108p 0 217.028p 0 217.029p 10000.0u 217.03p 0 221.285p 0 221.286p 10000.0u 221.287p 0 225.974p 0 225.975p 10000.0u 225.976p 0 239.084p 0 239.085p 10000.0u 239.086p 0 247.535p 0 247.536p 10000.0u 247.537p 0 260.117p 0 260.118p 10000.0u 260.119p 0 285.086p 0 285.087p 10000.0u 285.088p 0 288.617p 0 288.618p 10000.0u 288.619p 0 294.962p 0 294.963p 10000.0u 294.964p 0 302.978p 0 302.979p 10000.0u 302.98p 0 311.639p 0 311.64p 10000.0u 311.641p 0 322.475p 0 322.476p 10000.0u 322.477p 0 343.67p 0 343.671p 10000.0u 343.672p 0 344.573p 0 344.574p 10000.0u 344.575p 0 351.356p 0 351.357p 10000.0u 351.358p 0 353.045p 0 353.046p 10000.0u 353.047p 0 354.152p 0 354.153p 10000.0u 354.154p 0 357.113p 0 357.114p 10000.0u 357.115p 0 366.503p 0 366.504p 10000.0u 366.505p 0 375.041p 0 375.042p 10000.0u 375.043p 0 409.886p 0 409.887p 10000.0u 409.888p 0 411.548p 0 411.549p 10000.0u 411.55p 0 436.094p 0 436.095p 10000.0u 436.096p 0 442.7p 0 442.701p 10000.0u 442.702p 0 451.973p 0 451.974p 10000.0u 451.975p 0 452.924p 0 452.925p 10000.0u 452.926p 0 462.596p 0 462.597p 10000.0u 462.598p 0 476.246p 0 476.247p 10000.0u 476.248p 0 476.981p 0 476.982p 10000.0u 476.983p 0 478.916p 0 478.917p 10000.0u 478.918p 0 484.742p 0 484.743p 10000.0u 484.744p 0 485.576p 0 485.577p 10000.0u 485.578p 0 521.18p 0 521.181p 10000.0u 521.182p 0 526.838p 0 526.839p 10000.0u 526.84p 0 540.695p 0 540.696p 10000.0u 540.697p 0 541.133p 0 541.134p 10000.0u 541.135p 0 552.422p 0 552.423p 10000.0u 552.424p 0 556.073p 0 556.074p 10000.0u 556.075p 0 556.778p 0 556.779p 10000.0u 556.78p 0 573.926p 0 573.927p 10000.0u 573.928p 0 574.04p 0 574.041p 10000.0u 574.042p 0 576.839p 0 576.84p 10000.0u 576.841p 0 595.742p 0 595.743p 10000.0u 595.744p 0 596.681p 0 596.682p 10000.0u 596.683p 0 616.961p 0 616.962p 10000.0u 616.963p 0 623.162p 0 623.163p 10000.0u 623.164p 0 630.416p 0 630.417p 10000.0u 630.418p 0 654.518p 0 654.519p 10000.0u 654.52p 0 662.795p 0 662.796p 10000.0u 662.797p 0 677.729p 0 677.73p 10000.0u 677.731p 0 683.297p 0 683.298p 10000.0u 683.299p 0 690.485p 0 690.486p 10000.0u 690.487p 0 711.458p 0 711.459p 10000.0u 711.46p 0 716.729p 0 716.73p 10000.0u 716.731p 0 765.959p 0 765.96p 10000.0u 765.961p 0 782.879p 0 782.88p 10000.0u 782.881p 0 784.991p 0 784.992p 10000.0u 784.993p 0 804.302p 0 804.303p 10000.0u 804.304p 0 807.671p 0 807.672p 10000.0u 807.673p 0 809.153p 0 809.154p 10000.0u 809.155p 0 810.239p 0 810.24p 10000.0u 810.241p 0 824.246p 0 824.247p 10000.0u 824.248p 0 838.589p 0 838.59p 10000.0u 838.591p 0 862.451p 0 862.452p 10000.0u 862.453p 0 879.953p 0 879.954p 10000.0u 879.955p 0 881.102p 0 881.103p 10000.0u 881.104p 0 887.861p 0 887.862p 10000.0u 887.863p 0 900.296p 0 900.297p 10000.0u 900.298p 0 900.677p 0 900.678p 10000.0u 900.679p 0 904.787p 0 904.788p 10000.0u 904.789p 0 906.17p 0 906.171p 10000.0u 906.172p 0 927.365p 0 927.366p 10000.0u 927.367p 0 954.122p 0 954.123p 10000.0u 954.124p 0 961.331p 0 961.332p 10000.0u 961.333p 0 979.196p 0 979.197p 10000.0u 979.198p 0 982.478p 0 982.479p 10000.0u 982.48p 0 997.316p 0 997.317p 10000.0u 997.318p 0)
IIN79 0 80 pwl(0 0 21.596p 0 21.597p 10000.0u 21.598p 0 25.304p 0 25.305p 10000.0u 25.306p 0 33.536p 0 33.537p 10000.0u 33.538p 0 37.514p 0 37.515p 10000.0u 37.516p 0 38.3p 0 38.301p 10000.0u 38.302p 0 44.435p 0 44.436p 10000.0u 44.437p 0 47.315p 0 47.316p 10000.0u 47.317p 0 75.158p 0 75.159p 10000.0u 75.16p 0 75.425p 0 75.426p 10000.0u 75.427p 0 114.05p 0 114.051p 10000.0u 114.052p 0 136.703p 0 136.704p 10000.0u 136.705p 0 172.232p 0 172.233p 10000.0u 172.234p 0 192.257p 0 192.258p 10000.0u 192.259p 0 199.799p 0 199.8p 10000.0u 199.801p 0 201.35p 0 201.351p 10000.0u 201.352p 0 206.798p 0 206.799p 10000.0u 206.8p 0 222.989p 0 222.99p 10000.0u 222.991p 0 243.281p 0 243.282p 10000.0u 243.283p 0 292.928p 0 292.929p 10000.0u 292.93p 0 332.921p 0 332.922p 10000.0u 332.923p 0 352.724p 0 352.725p 10000.0u 352.726p 0 362.618p 0 362.619p 10000.0u 362.62p 0 367.211p 0 367.212p 10000.0u 367.213p 0 391.712p 0 391.713p 10000.0u 391.714p 0 409.88p 0 409.881p 10000.0u 409.882p 0 410.591p 0 410.592p 10000.0u 410.593p 0 429.083p 0 429.084p 10000.0u 429.085p 0 434.411p 0 434.412p 10000.0u 434.413p 0 434.948p 0 434.949p 10000.0u 434.95p 0 451.724p 0 451.725p 10000.0u 451.726p 0 468.386p 0 468.387p 10000.0u 468.388p 0 471.233p 0 471.234p 10000.0u 471.235p 0 477.824p 0 477.825p 10000.0u 477.826p 0 479.054p 0 479.055p 10000.0u 479.056p 0 490.469p 0 490.47p 10000.0u 490.471p 0 503.087p 0 503.088p 10000.0u 503.089p 0 504.686p 0 504.687p 10000.0u 504.688p 0 521.294p 0 521.295p 10000.0u 521.296p 0 535.556p 0 535.557p 10000.0u 535.558p 0 538.22p 0 538.221p 10000.0u 538.222p 0 566.732p 0 566.733p 10000.0u 566.734p 0 579.014p 0 579.015p 10000.0u 579.016p 0 579.779p 0 579.78p 10000.0u 579.781p 0 584.999p 0 585.0p 10000.0u 585.001p 0 591.782p 0 591.783p 10000.0u 591.784p 0 595.067p 0 595.068p 10000.0u 595.069p 0 613.91p 0 613.911p 10000.0u 613.912p 0 617.885p 0 617.886p 10000.0u 617.887p 0 629.27p 0 629.271p 10000.0u 629.272p 0 642.749p 0 642.75p 10000.0u 642.751p 0 643.166p 0 643.167p 10000.0u 643.168p 0 646.808p 0 646.809p 10000.0u 646.81p 0 654.875p 0 654.876p 10000.0u 654.877p 0 672.515p 0 672.516p 10000.0u 672.517p 0 682.889p 0 682.89p 10000.0u 682.891p 0 685.754p 0 685.755p 10000.0u 685.756p 0 686.879p 0 686.88p 10000.0u 686.881p 0 693.578p 0 693.579p 10000.0u 693.58p 0 701.105p 0 701.106p 10000.0u 701.107p 0 702.989p 0 702.99p 10000.0u 702.991p 0 704.573p 0 704.574p 10000.0u 704.575p 0 704.804p 0 704.805p 10000.0u 704.806p 0 719.777p 0 719.778p 10000.0u 719.779p 0 720.944p 0 720.945p 10000.0u 720.946p 0 723.578p 0 723.579p 10000.0u 723.58p 0 723.626p 0 723.627p 10000.0u 723.628p 0 744.908p 0 744.909p 10000.0u 744.91p 0 746.021p 0 746.022p 10000.0u 746.023p 0 752.186p 0 752.187p 10000.0u 752.188p 0 753.269p 0 753.27p 10000.0u 753.271p 0 776.423p 0 776.424p 10000.0u 776.425p 0 783.926p 0 783.927p 10000.0u 783.928p 0 795.905p 0 795.906p 10000.0u 795.907p 0 817.712p 0 817.713p 10000.0u 817.714p 0 833.39p 0 833.391p 10000.0u 833.392p 0 839.735p 0 839.736p 10000.0u 839.737p 0 852.098p 0 852.099p 10000.0u 852.1p 0 857.408p 0 857.409p 10000.0u 857.41p 0 869.438p 0 869.439p 10000.0u 869.44p 0 875.165p 0 875.166p 10000.0u 875.167p 0 876.14p 0 876.141p 10000.0u 876.142p 0 894.983p 0 894.984p 10000.0u 894.985p 0 929.894p 0 929.895p 10000.0u 929.896p 0 929.933p 0 929.934p 10000.0u 929.935p 0 937.694p 0 937.695p 10000.0u 937.696p 0 942.143p 0 942.144p 10000.0u 942.145p 0 947.702p 0 947.703p 10000.0u 947.704p 0 949.643p 0 949.644p 10000.0u 949.645p 0 953.843p 0 953.844p 10000.0u 953.845p 0 970.061p 0 970.062p 10000.0u 970.063p 0 993.038p 0 993.039p 10000.0u 993.04p 0 993.887p 0 993.888p 10000.0u 993.889p 0)
IIN80 0 81 pwl(0 0 6.851p 0 6.852p 10000.0u 6.853p 0 7.172p 0 7.173p 10000.0u 7.174p 0 21.743p 0 21.744p 10000.0u 21.745p 0 26.78p 0 26.781p 10000.0u 26.782p 0 29.945p 0 29.946p 10000.0u 29.947p 0 56.669p 0 56.67p 10000.0u 56.671p 0 64.511p 0 64.512p 10000.0u 64.513p 0 76.931p 0 76.932p 10000.0u 76.933p 0 81.314p 0 81.315p 10000.0u 81.316p 0 90.173p 0 90.174p 10000.0u 90.175p 0 102.71p 0 102.711p 10000.0u 102.712p 0 127.973p 0 127.974p 10000.0u 127.975p 0 139.574p 0 139.575p 10000.0u 139.576p 0 153.938p 0 153.939p 10000.0u 153.94p 0 155.531p 0 155.532p 10000.0u 155.533p 0 161.903p 0 161.904p 10000.0u 161.905p 0 166.055p 0 166.056p 10000.0u 166.057p 0 167.093p 0 167.094p 10000.0u 167.095p 0 169.901p 0 169.902p 10000.0u 169.903p 0 171.509p 0 171.51p 10000.0u 171.511p 0 173.063p 0 173.064p 10000.0u 173.065p 0 183.188p 0 183.189p 10000.0u 183.19p 0 183.761p 0 183.762p 10000.0u 183.763p 0 185.066p 0 185.067p 10000.0u 185.068p 0 190.802p 0 190.803p 10000.0u 190.804p 0 198.866p 0 198.867p 10000.0u 198.868p 0 201.326p 0 201.327p 10000.0u 201.328p 0 203.87p 0 203.871p 10000.0u 203.872p 0 231.722p 0 231.723p 10000.0u 231.724p 0 234.644p 0 234.645p 10000.0u 234.646p 0 247.199p 0 247.2p 10000.0u 247.201p 0 247.898p 0 247.899p 10000.0u 247.9p 0 252.947p 0 252.948p 10000.0u 252.949p 0 263.819p 0 263.82p 10000.0u 263.821p 0 271.193p 0 271.194p 10000.0u 271.195p 0 274.904p 0 274.905p 10000.0u 274.906p 0 277.004p 0 277.005p 10000.0u 277.006p 0 283.304p 0 283.305p 10000.0u 283.306p 0 303.269p 0 303.27p 10000.0u 303.271p 0 306.377p 0 306.378p 10000.0u 306.379p 0 342.635p 0 342.636p 10000.0u 342.637p 0 345.149p 0 345.15p 10000.0u 345.151p 0 351.305p 0 351.306p 10000.0u 351.307p 0 354.734p 0 354.735p 10000.0u 354.736p 0 356.012p 0 356.013p 10000.0u 356.014p 0 362.408p 0 362.409p 10000.0u 362.41p 0 363.758p 0 363.759p 10000.0u 363.76p 0 370.145p 0 370.146p 10000.0u 370.147p 0 390.245p 0 390.246p 10000.0u 390.247p 0 397.964p 0 397.965p 10000.0u 397.966p 0 405.734p 0 405.735p 10000.0u 405.736p 0 414.038p 0 414.039p 10000.0u 414.04p 0 453.917p 0 453.918p 10000.0u 453.919p 0 455.084p 0 455.085p 10000.0u 455.086p 0 463.142p 0 463.143p 10000.0u 463.144p 0 479.696p 0 479.697p 10000.0u 479.698p 0 484.886p 0 484.887p 10000.0u 484.888p 0 494.339p 0 494.34p 10000.0u 494.341p 0 495.875p 0 495.876p 10000.0u 495.877p 0 518.102p 0 518.103p 10000.0u 518.104p 0 533.006p 0 533.007p 10000.0u 533.008p 0 538.313p 0 538.314p 10000.0u 538.315p 0 556.355p 0 556.356p 10000.0u 556.357p 0 563.822p 0 563.823p 10000.0u 563.824p 0 565.874p 0 565.875p 10000.0u 565.876p 0 571.067p 0 571.068p 10000.0u 571.069p 0 580.661p 0 580.662p 10000.0u 580.663p 0 581.819p 0 581.82p 10000.0u 581.821p 0 596.402p 0 596.403p 10000.0u 596.404p 0 615.341p 0 615.342p 10000.0u 615.343p 0 639.617p 0 639.618p 10000.0u 639.619p 0 642.578p 0 642.579p 10000.0u 642.58p 0 643.379p 0 643.38p 10000.0u 643.381p 0 673.094p 0 673.095p 10000.0u 673.096p 0 674.411p 0 674.412p 10000.0u 674.413p 0 692.225p 0 692.226p 10000.0u 692.227p 0 700.208p 0 700.209p 10000.0u 700.21p 0 700.988p 0 700.989p 10000.0u 700.99p 0 704.255p 0 704.256p 10000.0u 704.257p 0 766.205p 0 766.206p 10000.0u 766.207p 0 774.806p 0 774.807p 10000.0u 774.808p 0 777.053p 0 777.054p 10000.0u 777.055p 0 795.926p 0 795.927p 10000.0u 795.928p 0 817.88p 0 817.881p 10000.0u 817.882p 0 825.311p 0 825.312p 10000.0u 825.313p 0 827.03p 0 827.031p 10000.0u 827.032p 0 829.082p 0 829.083p 10000.0u 829.084p 0 835.019p 0 835.02p 10000.0u 835.021p 0 836.552p 0 836.553p 10000.0u 836.554p 0 847.325p 0 847.326p 10000.0u 847.327p 0 851.972p 0 851.973p 10000.0u 851.974p 0 854.519p 0 854.52p 10000.0u 854.521p 0 862.589p 0 862.59p 10000.0u 862.591p 0 896.21p 0 896.211p 10000.0u 896.212p 0 896.591p 0 896.592p 10000.0u 896.593p 0 901.928p 0 901.929p 10000.0u 901.93p 0 902.195p 0 902.196p 10000.0u 902.197p 0 909.755p 0 909.756p 10000.0u 909.757p 0 921.161p 0 921.162p 10000.0u 921.163p 0 926.432p 0 926.433p 10000.0u 926.434p 0 927.875p 0 927.876p 10000.0u 927.877p 0 950.189p 0 950.19p 10000.0u 950.191p 0 975.02p 0 975.021p 10000.0u 975.022p 0 999.515p 0 999.516p 10000.0u 999.517p 0)
IIN81 0 82 pwl(0 0 34.502p 0 34.503p 10000.0u 34.504p 0 35.606p 0 35.607p 10000.0u 35.608p 0 48.116p 0 48.117p 10000.0u 48.118p 0 58.979p 0 58.98p 10000.0u 58.981p 0 73.133p 0 73.134p 10000.0u 73.135p 0 81.701p 0 81.702p 10000.0u 81.703p 0 94.43p 0 94.431p 10000.0u 94.432p 0 97.169p 0 97.17p 10000.0u 97.171p 0 119.396p 0 119.397p 10000.0u 119.398p 0 133.349p 0 133.35p 10000.0u 133.351p 0 143.42p 0 143.421p 10000.0u 143.422p 0 143.753p 0 143.754p 10000.0u 143.755p 0 146.009p 0 146.01p 10000.0u 146.011p 0 189.017p 0 189.018p 10000.0u 189.019p 0 203.714p 0 203.715p 10000.0u 203.716p 0 207.92p 0 207.921p 10000.0u 207.922p 0 217.514p 0 217.515p 10000.0u 217.516p 0 220.076p 0 220.077p 10000.0u 220.078p 0 230.363p 0 230.364p 10000.0u 230.365p 0 252.578p 0 252.579p 10000.0u 252.58p 0 254.963p 0 254.964p 10000.0u 254.965p 0 266.006p 0 266.007p 10000.0u 266.008p 0 270.035p 0 270.036p 10000.0u 270.037p 0 273.218p 0 273.219p 10000.0u 273.22p 0 308.645p 0 308.646p 10000.0u 308.647p 0 308.918p 0 308.919p 10000.0u 308.92p 0 311.255p 0 311.256p 10000.0u 311.257p 0 312.011p 0 312.012p 10000.0u 312.013p 0 321.671p 0 321.672p 10000.0u 321.673p 0 326.408p 0 326.409p 10000.0u 326.41p 0 347.069p 0 347.07p 10000.0u 347.071p 0 349.445p 0 349.446p 10000.0u 349.447p 0 351.02p 0 351.021p 10000.0u 351.022p 0 360.089p 0 360.09p 10000.0u 360.091p 0 360.779p 0 360.78p 10000.0u 360.781p 0 362.318p 0 362.319p 10000.0u 362.32p 0 379.478p 0 379.479p 10000.0u 379.48p 0 380.339p 0 380.34p 10000.0u 380.341p 0 382.91p 0 382.911p 10000.0u 382.912p 0 383.375p 0 383.376p 10000.0u 383.377p 0 414.02p 0 414.021p 10000.0u 414.022p 0 414.104p 0 414.105p 10000.0u 414.106p 0 423.857p 0 423.858p 10000.0u 423.859p 0 429.977p 0 429.978p 10000.0u 429.979p 0 438.398p 0 438.399p 10000.0u 438.4p 0 462.902p 0 462.903p 10000.0u 462.904p 0 466.451p 0 466.452p 10000.0u 466.453p 0 471.593p 0 471.594p 10000.0u 471.595p 0 473.072p 0 473.073p 10000.0u 473.074p 0 476.99p 0 476.991p 10000.0u 476.992p 0 477.614p 0 477.615p 10000.0u 477.616p 0 481.961p 0 481.962p 10000.0u 481.963p 0 484.79p 0 484.791p 10000.0u 484.792p 0 496.859p 0 496.86p 10000.0u 496.861p 0 500.552p 0 500.553p 10000.0u 500.554p 0 515.6p 0 515.601p 10000.0u 515.602p 0 518.375p 0 518.376p 10000.0u 518.377p 0 544.328p 0 544.329p 10000.0u 544.33p 0 570.791p 0 570.792p 10000.0u 570.793p 0 583.376p 0 583.377p 10000.0u 583.378p 0 600.914p 0 600.915p 10000.0u 600.916p 0 612.572p 0 612.573p 10000.0u 612.574p 0 613.517p 0 613.518p 10000.0u 613.519p 0 636.53p 0 636.531p 10000.0u 636.532p 0 639.074p 0 639.075p 10000.0u 639.076p 0 647.417p 0 647.418p 10000.0u 647.419p 0 648.917p 0 648.918p 10000.0u 648.919p 0 662.501p 0 662.502p 10000.0u 662.503p 0 667.613p 0 667.614p 10000.0u 667.615p 0 668.408p 0 668.409p 10000.0u 668.41p 0 670.469p 0 670.47p 10000.0u 670.471p 0 675.386p 0 675.387p 10000.0u 675.388p 0 682.172p 0 682.173p 10000.0u 682.174p 0 695.804p 0 695.805p 10000.0u 695.806p 0 697.01p 0 697.011p 10000.0u 697.012p 0 700.589p 0 700.59p 10000.0u 700.591p 0 703.415p 0 703.416p 10000.0u 703.417p 0 718.52p 0 718.521p 10000.0u 718.522p 0 730.25p 0 730.251p 10000.0u 730.252p 0 735.32p 0 735.321p 10000.0u 735.322p 0 739.811p 0 739.812p 10000.0u 739.813p 0 741.074p 0 741.075p 10000.0u 741.076p 0 778.247p 0 778.248p 10000.0u 778.249p 0 790.394p 0 790.395p 10000.0u 790.396p 0 792.839p 0 792.84p 10000.0u 792.841p 0 801.365p 0 801.366p 10000.0u 801.367p 0 820.739p 0 820.74p 10000.0u 820.741p 0 821.633p 0 821.634p 10000.0u 821.635p 0 831.95p 0 831.951p 10000.0u 831.952p 0 832.037p 0 832.038p 10000.0u 832.039p 0 833.588p 0 833.589p 10000.0u 833.59p 0 838.124p 0 838.125p 10000.0u 838.126p 0 840.434p 0 840.435p 10000.0u 840.436p 0 843.398p 0 843.399p 10000.0u 843.4p 0 870.089p 0 870.09p 10000.0u 870.091p 0 877.445p 0 877.446p 10000.0u 877.447p 0 882.119p 0 882.12p 10000.0u 882.121p 0 890.294p 0 890.295p 10000.0u 890.296p 0 900.719p 0 900.72p 10000.0u 900.721p 0 905.906p 0 905.907p 10000.0u 905.908p 0 924.896p 0 924.897p 10000.0u 924.898p 0 933.803p 0 933.804p 10000.0u 933.805p 0 934.952p 0 934.953p 10000.0u 934.954p 0 948.011p 0 948.012p 10000.0u 948.013p 0 954.02p 0 954.021p 10000.0u 954.022p 0 987.926p 0 987.927p 10000.0u 987.928p 0)
IIN82 0 83 pwl(0 0 6.404p 0 6.405p 10000.0u 6.406p 0 9.014p 0 9.015p 10000.0u 9.016p 0 28.376p 0 28.377p 10000.0u 28.378p 0 50.312p 0 50.313p 10000.0u 50.314p 0 56.828p 0 56.829p 10000.0u 56.83p 0 81.116p 0 81.117p 10000.0u 81.118p 0 90.506p 0 90.507p 10000.0u 90.508p 0 90.782p 0 90.783p 10000.0u 90.784p 0 102.662p 0 102.663p 10000.0u 102.664p 0 119.891p 0 119.892p 10000.0u 119.893p 0 121.271p 0 121.272p 10000.0u 121.273p 0 123.035p 0 123.036p 10000.0u 123.037p 0 139.496p 0 139.497p 10000.0u 139.498p 0 139.544p 0 139.545p 10000.0u 139.546p 0 142.61p 0 142.611p 10000.0u 142.612p 0 145.679p 0 145.68p 10000.0u 145.681p 0 153.563p 0 153.564p 10000.0u 153.565p 0 155.588p 0 155.589p 10000.0u 155.59p 0 162.104p 0 162.105p 10000.0u 162.106p 0 198.467p 0 198.468p 10000.0u 198.469p 0 201.017p 0 201.018p 10000.0u 201.019p 0 209.621p 0 209.622p 10000.0u 209.623p 0 224.06p 0 224.061p 10000.0u 224.062p 0 225.248p 0 225.249p 10000.0u 225.25p 0 254.816p 0 254.817p 10000.0u 254.818p 0 268.079p 0 268.08p 10000.0u 268.081p 0 280.757p 0 280.758p 10000.0u 280.759p 0 289.211p 0 289.212p 10000.0u 289.213p 0 294.584p 0 294.585p 10000.0u 294.586p 0 306.62p 0 306.621p 10000.0u 306.622p 0 314.498p 0 314.499p 10000.0u 314.5p 0 333.209p 0 333.21p 10000.0u 333.211p 0 341.714p 0 341.715p 10000.0u 341.716p 0 344.363p 0 344.364p 10000.0u 344.365p 0 349.157p 0 349.158p 10000.0u 349.159p 0 354.281p 0 354.282p 10000.0u 354.283p 0 359.219p 0 359.22p 10000.0u 359.221p 0 370.883p 0 370.884p 10000.0u 370.885p 0 385.538p 0 385.539p 10000.0u 385.54p 0 386.384p 0 386.385p 10000.0u 386.386p 0 417.515p 0 417.516p 10000.0u 417.517p 0 431.318p 0 431.319p 10000.0u 431.32p 0 432.287p 0 432.288p 10000.0u 432.289p 0 434.297p 0 434.298p 10000.0u 434.299p 0 439.004p 0 439.005p 10000.0u 439.006p 0 461.081p 0 461.082p 10000.0u 461.083p 0 466.244p 0 466.245p 10000.0u 466.246p 0 496.589p 0 496.59p 10000.0u 496.591p 0 500.987p 0 500.988p 10000.0u 500.989p 0 516.641p 0 516.642p 10000.0u 516.643p 0 526.94p 0 526.941p 10000.0u 526.942p 0 527.429p 0 527.43p 10000.0u 527.431p 0 542.87p 0 542.871p 10000.0u 542.872p 0 568.442p 0 568.443p 10000.0u 568.444p 0 574.796p 0 574.797p 10000.0u 574.798p 0 611.243p 0 611.244p 10000.0u 611.245p 0 614.609p 0 614.61p 10000.0u 614.611p 0 638.876p 0 638.877p 10000.0u 638.878p 0 650.639p 0 650.64p 10000.0u 650.641p 0 667.676p 0 667.677p 10000.0u 667.678p 0 667.931p 0 667.932p 10000.0u 667.933p 0 674.408p 0 674.409p 10000.0u 674.41p 0 677.042p 0 677.043p 10000.0u 677.044p 0 680.339p 0 680.34p 10000.0u 680.341p 0 682.463p 0 682.464p 10000.0u 682.465p 0 689.06p 0 689.061p 10000.0u 689.062p 0 696.671p 0 696.672p 10000.0u 696.673p 0 716.558p 0 716.559p 10000.0u 716.56p 0 725.285p 0 725.286p 10000.0u 725.287p 0 728.384p 0 728.385p 10000.0u 728.386p 0 728.756p 0 728.757p 10000.0u 728.758p 0 736.295p 0 736.296p 10000.0u 736.297p 0 740.735p 0 740.736p 10000.0u 740.737p 0 742.031p 0 742.032p 10000.0u 742.033p 0 758.129p 0 758.13p 10000.0u 758.131p 0 784.502p 0 784.503p 10000.0u 784.504p 0 813.026p 0 813.027p 10000.0u 813.028p 0 825.476p 0 825.477p 10000.0u 825.478p 0 831.629p 0 831.63p 10000.0u 831.631p 0 848.897p 0 848.898p 10000.0u 848.899p 0 858.599p 0 858.6p 10000.0u 858.601p 0 871.7p 0 871.701p 10000.0u 871.702p 0 873.653p 0 873.654p 10000.0u 873.655p 0 878.651p 0 878.652p 10000.0u 878.653p 0 880.388p 0 880.389p 10000.0u 880.39p 0 915.959p 0 915.96p 10000.0u 915.961p 0 917.72p 0 917.721p 10000.0u 917.722p 0 949.634p 0 949.635p 10000.0u 949.636p 0 988.007p 0 988.008p 10000.0u 988.009p 0 988.208p 0 988.209p 10000.0u 988.21p 0 999.188p 0 999.189p 10000.0u 999.19p 0)
IIN83 0 84 pwl(0 0 7.82p 0 7.821p 10000.0u 7.822p 0 12.662p 0 12.663p 10000.0u 12.664p 0 18.29p 0 18.291p 10000.0u 18.292p 0 32.969p 0 32.97p 10000.0u 32.971p 0 36.119p 0 36.12p 10000.0u 36.121p 0 40.88p 0 40.881p 10000.0u 40.882p 0 58.901p 0 58.902p 10000.0u 58.903p 0 63.983p 0 63.984p 10000.0u 63.985p 0 83.507p 0 83.508p 10000.0u 83.509p 0 93.473p 0 93.474p 10000.0u 93.475p 0 100.277p 0 100.278p 10000.0u 100.279p 0 101.735p 0 101.736p 10000.0u 101.737p 0 120.332p 0 120.333p 10000.0u 120.334p 0 127.922p 0 127.923p 10000.0u 127.924p 0 128.528p 0 128.529p 10000.0u 128.53p 0 138.95p 0 138.951p 10000.0u 138.952p 0 147.737p 0 147.738p 10000.0u 147.739p 0 169.34p 0 169.341p 10000.0u 169.342p 0 191.159p 0 191.16p 10000.0u 191.161p 0 191.39p 0 191.391p 10000.0u 191.392p 0 211.391p 0 211.392p 10000.0u 211.393p 0 215.528p 0 215.529p 10000.0u 215.53p 0 220.682p 0 220.683p 10000.0u 220.684p 0 263.837p 0 263.838p 10000.0u 263.839p 0 270.08p 0 270.081p 10000.0u 270.082p 0 274.643p 0 274.644p 10000.0u 274.645p 0 274.958p 0 274.959p 10000.0u 274.96p 0 290.3p 0 290.301p 10000.0u 290.302p 0 290.696p 0 290.697p 10000.0u 290.698p 0 295.949p 0 295.95p 10000.0u 295.951p 0 300.233p 0 300.234p 10000.0u 300.235p 0 303.287p 0 303.288p 10000.0u 303.289p 0 303.839p 0 303.84p 10000.0u 303.841p 0 317.717p 0 317.718p 10000.0u 317.719p 0 318.278p 0 318.279p 10000.0u 318.28p 0 319.976p 0 319.977p 10000.0u 319.978p 0 329.231p 0 329.232p 10000.0u 329.233p 0 329.315p 0 329.316p 10000.0u 329.317p 0 335.582p 0 335.583p 10000.0u 335.584p 0 341.18p 0 341.181p 10000.0u 341.182p 0 342.149p 0 342.15p 10000.0u 342.151p 0 354.527p 0 354.528p 10000.0u 354.529p 0 362.342p 0 362.343p 10000.0u 362.344p 0 365.429p 0 365.43p 10000.0u 365.431p 0 391.217p 0 391.218p 10000.0u 391.219p 0 396.704p 0 396.705p 10000.0u 396.706p 0 399.266p 0 399.267p 10000.0u 399.268p 0 408.269p 0 408.27p 10000.0u 408.271p 0 435.212p 0 435.213p 10000.0u 435.214p 0 441.128p 0 441.129p 10000.0u 441.13p 0 443.192p 0 443.193p 10000.0u 443.194p 0 474.665p 0 474.666p 10000.0u 474.667p 0 482.009p 0 482.01p 10000.0u 482.011p 0 494.822p 0 494.823p 10000.0u 494.824p 0 497.291p 0 497.292p 10000.0u 497.293p 0 498.743p 0 498.744p 10000.0u 498.745p 0 501.251p 0 501.252p 10000.0u 501.253p 0 502.721p 0 502.722p 10000.0u 502.723p 0 514.514p 0 514.515p 10000.0u 514.516p 0 524.447p 0 524.448p 10000.0u 524.449p 0 533.879p 0 533.88p 10000.0u 533.881p 0 543.845p 0 543.846p 10000.0u 543.847p 0 547.133p 0 547.134p 10000.0u 547.135p 0 550.055p 0 550.056p 10000.0u 550.057p 0 556.508p 0 556.509p 10000.0u 556.51p 0 559.274p 0 559.275p 10000.0u 559.276p 0 561.035p 0 561.036p 10000.0u 561.037p 0 565.961p 0 565.962p 10000.0u 565.963p 0 578.723p 0 578.724p 10000.0u 578.725p 0 617.513p 0 617.514p 10000.0u 617.515p 0 617.6p 0 617.601p 10000.0u 617.602p 0 623.996p 0 623.997p 10000.0u 623.998p 0 624.542p 0 624.543p 10000.0u 624.544p 0 636.092p 0 636.093p 10000.0u 636.094p 0 644.054p 0 644.055p 10000.0u 644.056p 0 653.462p 0 653.463p 10000.0u 653.464p 0 678.035p 0 678.036p 10000.0u 678.037p 0 696.041p 0 696.042p 10000.0u 696.043p 0 708.884p 0 708.885p 10000.0u 708.886p 0 729.788p 0 729.789p 10000.0u 729.79p 0 738.551p 0 738.552p 10000.0u 738.553p 0 739.943p 0 739.944p 10000.0u 739.945p 0 742.604p 0 742.605p 10000.0u 742.606p 0 753.029p 0 753.03p 10000.0u 753.031p 0 760.22p 0 760.221p 10000.0u 760.222p 0 776.009p 0 776.01p 10000.0u 776.011p 0 783.485p 0 783.486p 10000.0u 783.487p 0 790.382p 0 790.383p 10000.0u 790.384p 0 801.041p 0 801.042p 10000.0u 801.043p 0 809.45p 0 809.451p 10000.0u 809.452p 0 816.656p 0 816.657p 10000.0u 816.658p 0 817.304p 0 817.305p 10000.0u 817.306p 0 826.205p 0 826.206p 10000.0u 826.207p 0 850.892p 0 850.893p 10000.0u 850.894p 0 851.903p 0 851.904p 10000.0u 851.905p 0 862.106p 0 862.107p 10000.0u 862.108p 0 866.924p 0 866.925p 10000.0u 866.926p 0 878.354p 0 878.355p 10000.0u 878.356p 0 884.741p 0 884.742p 10000.0u 884.743p 0 904.154p 0 904.155p 10000.0u 904.156p 0 905.621p 0 905.622p 10000.0u 905.623p 0 917.675p 0 917.676p 10000.0u 917.677p 0 942.599p 0 942.6p 10000.0u 942.601p 0 965.174p 0 965.175p 10000.0u 965.176p 0 968.189p 0 968.19p 10000.0u 968.191p 0 980.627p 0 980.628p 10000.0u 980.629p 0)
IIN84 0 85 pwl(0 0 1.052p 0 1.053p 10000.0u 1.054p 0 74.18p 0 74.181p 10000.0u 74.182p 0 85.262p 0 85.263p 10000.0u 85.264p 0 86.774p 0 86.775p 10000.0u 86.776p 0 100.682p 0 100.683p 10000.0u 100.684p 0 118.391p 0 118.392p 10000.0u 118.393p 0 147.935p 0 147.936p 10000.0u 147.937p 0 161.804p 0 161.805p 10000.0u 161.806p 0 166.448p 0 166.449p 10000.0u 166.45p 0 167.864p 0 167.865p 10000.0u 167.866p 0 185.174p 0 185.175p 10000.0u 185.176p 0 202.511p 0 202.512p 10000.0u 202.513p 0 211.007p 0 211.008p 10000.0u 211.009p 0 212.762p 0 212.763p 10000.0u 212.764p 0 217.607p 0 217.608p 10000.0u 217.609p 0 218.798p 0 218.799p 10000.0u 218.8p 0 240.029p 0 240.03p 10000.0u 240.031p 0 241.637p 0 241.638p 10000.0u 241.639p 0 241.778p 0 241.779p 10000.0u 241.78p 0 245.63p 0 245.631p 10000.0u 245.632p 0 246.23p 0 246.231p 10000.0u 246.232p 0 253.613p 0 253.614p 10000.0u 253.615p 0 266.612p 0 266.613p 10000.0u 266.614p 0 272.114p 0 272.115p 10000.0u 272.116p 0 274.961p 0 274.962p 10000.0u 274.963p 0 281.756p 0 281.757p 10000.0u 281.758p 0 281.771p 0 281.772p 10000.0u 281.773p 0 293.423p 0 293.424p 10000.0u 293.425p 0 298.856p 0 298.857p 10000.0u 298.858p 0 301.076p 0 301.077p 10000.0u 301.078p 0 314.51p 0 314.511p 10000.0u 314.512p 0 336.545p 0 336.546p 10000.0u 336.547p 0 338.081p 0 338.082p 10000.0u 338.083p 0 342.401p 0 342.402p 10000.0u 342.403p 0 350.735p 0 350.736p 10000.0u 350.737p 0 352.199p 0 352.2p 10000.0u 352.201p 0 364.064p 0 364.065p 10000.0u 364.066p 0 371.789p 0 371.79p 10000.0u 371.791p 0 377.498p 0 377.499p 10000.0u 377.5p 0 418.295p 0 418.296p 10000.0u 418.297p 0 431.33p 0 431.331p 10000.0u 431.332p 0 455.36p 0 455.361p 10000.0u 455.362p 0 467.225p 0 467.226p 10000.0u 467.227p 0 471.257p 0 471.258p 10000.0u 471.259p 0 477.815p 0 477.816p 10000.0u 477.817p 0 496.955p 0 496.956p 10000.0u 496.957p 0 497.99p 0 497.991p 10000.0u 497.992p 0 525.548p 0 525.549p 10000.0u 525.55p 0 552.701p 0 552.702p 10000.0u 552.703p 0 553.238p 0 553.239p 10000.0u 553.24p 0 555.866p 0 555.867p 10000.0u 555.868p 0 564.782p 0 564.783p 10000.0u 564.784p 0 565.502p 0 565.503p 10000.0u 565.504p 0 572.798p 0 572.799p 10000.0u 572.8p 0 577.769p 0 577.77p 10000.0u 577.771p 0 599.42p 0 599.421p 10000.0u 599.422p 0 609.335p 0 609.336p 10000.0u 609.337p 0 613.808p 0 613.809p 10000.0u 613.81p 0 617.825p 0 617.826p 10000.0u 617.827p 0 618.308p 0 618.309p 10000.0u 618.31p 0 639.542p 0 639.543p 10000.0u 639.544p 0 643.793p 0 643.794p 10000.0u 643.795p 0 671.441p 0 671.442p 10000.0u 671.443p 0 681.632p 0 681.633p 10000.0u 681.634p 0 683.399p 0 683.4p 10000.0u 683.401p 0 701.678p 0 701.679p 10000.0u 701.68p 0 728.594p 0 728.595p 10000.0u 728.596p 0 739.604p 0 739.605p 10000.0u 739.606p 0 740.888p 0 740.889p 10000.0u 740.89p 0 745.175p 0 745.176p 10000.0u 745.177p 0 810.245p 0 810.246p 10000.0u 810.247p 0 818.489p 0 818.49p 10000.0u 818.491p 0 821.474p 0 821.475p 10000.0u 821.476p 0 843.302p 0 843.303p 10000.0u 843.304p 0 851.318p 0 851.319p 10000.0u 851.32p 0 870.134p 0 870.135p 10000.0u 870.136p 0 892.025p 0 892.026p 10000.0u 892.027p 0 916.313p 0 916.314p 10000.0u 916.315p 0 919.841p 0 919.842p 10000.0u 919.843p 0 926.918p 0 926.919p 10000.0u 926.92p 0 953.474p 0 953.475p 10000.0u 953.476p 0 965.447p 0 965.448p 10000.0u 965.449p 0 969.44p 0 969.441p 10000.0u 969.442p 0 974.153p 0 974.154p 10000.0u 974.155p 0 978.167p 0 978.168p 10000.0u 978.169p 0 990.149p 0 990.15p 10000.0u 990.151p 0 994.667p 0 994.668p 10000.0u 994.669p 0)
IIN85 0 86 pwl(0 0 0.329p 0 0.33p 10000.0u 0.331p 0 4.724p 0 4.725p 10000.0u 4.726p 0 7.13p 0 7.131p 10000.0u 7.132p 0 10.133p 0 10.134p 10000.0u 10.135p 0 18.953p 0 18.954p 10000.0u 18.955p 0 25.604p 0 25.605p 10000.0u 25.606p 0 28.46p 0 28.461p 10000.0u 28.462p 0 30.884p 0 30.885p 10000.0u 30.886p 0 57.515p 0 57.516p 10000.0u 57.517p 0 57.686p 0 57.687p 10000.0u 57.688p 0 61.487p 0 61.488p 10000.0u 61.489p 0 81.428p 0 81.429p 10000.0u 81.43p 0 82.697p 0 82.698p 10000.0u 82.699p 0 84.23p 0 84.231p 10000.0u 84.232p 0 103.901p 0 103.902p 10000.0u 103.903p 0 108.356p 0 108.357p 10000.0u 108.358p 0 123.734p 0 123.735p 10000.0u 123.736p 0 125.312p 0 125.313p 10000.0u 125.314p 0 140.6p 0 140.601p 10000.0u 140.602p 0 149.774p 0 149.775p 10000.0u 149.776p 0 151.019p 0 151.02p 10000.0u 151.021p 0 155.657p 0 155.658p 10000.0u 155.659p 0 166.529p 0 166.53p 10000.0u 166.531p 0 210.377p 0 210.378p 10000.0u 210.379p 0 217.253p 0 217.254p 10000.0u 217.255p 0 220.874p 0 220.875p 10000.0u 220.876p 0 234.965p 0 234.966p 10000.0u 234.967p 0 237.659p 0 237.66p 10000.0u 237.661p 0 238.421p 0 238.422p 10000.0u 238.423p 0 239.132p 0 239.133p 10000.0u 239.134p 0 243.77p 0 243.771p 10000.0u 243.772p 0 244.355p 0 244.356p 10000.0u 244.357p 0 255.338p 0 255.339p 10000.0u 255.34p 0 263.552p 0 263.553p 10000.0u 263.554p 0 275.027p 0 275.028p 10000.0u 275.029p 0 281.171p 0 281.172p 10000.0u 281.173p 0 286.001p 0 286.002p 10000.0u 286.003p 0 299.939p 0 299.94p 10000.0u 299.941p 0 302.681p 0 302.682p 10000.0u 302.683p 0 305.789p 0 305.79p 10000.0u 305.791p 0 334.229p 0 334.23p 10000.0u 334.231p 0 343.601p 0 343.602p 10000.0u 343.603p 0 354.284p 0 354.285p 10000.0u 354.286p 0 379.307p 0 379.308p 10000.0u 379.309p 0 409.745p 0 409.746p 10000.0u 409.747p 0 409.952p 0 409.953p 10000.0u 409.954p 0 412.097p 0 412.098p 10000.0u 412.099p 0 427.97p 0 427.971p 10000.0u 427.972p 0 434.708p 0 434.709p 10000.0u 434.71p 0 460.565p 0 460.566p 10000.0u 460.567p 0 475.916p 0 475.917p 10000.0u 475.918p 0 478.673p 0 478.674p 10000.0u 478.675p 0 481.265p 0 481.266p 10000.0u 481.267p 0 511.694p 0 511.695p 10000.0u 511.696p 0 517.397p 0 517.398p 10000.0u 517.399p 0 523.724p 0 523.725p 10000.0u 523.726p 0 525.938p 0 525.939p 10000.0u 525.94p 0 531.038p 0 531.039p 10000.0u 531.04p 0 534.455p 0 534.456p 10000.0u 534.457p 0 543.506p 0 543.507p 10000.0u 543.508p 0 546.932p 0 546.933p 10000.0u 546.934p 0 565.34p 0 565.341p 10000.0u 565.342p 0 586.328p 0 586.329p 10000.0u 586.33p 0 597.806p 0 597.807p 10000.0u 597.808p 0 613.088p 0 613.089p 10000.0u 613.09p 0 614.546p 0 614.547p 10000.0u 614.548p 0 615.338p 0 615.339p 10000.0u 615.34p 0 628.55p 0 628.551p 10000.0u 628.552p 0 630.824p 0 630.825p 10000.0u 630.826p 0 641.867p 0 641.868p 10000.0u 641.869p 0 653.084p 0 653.085p 10000.0u 653.086p 0 656.168p 0 656.169p 10000.0u 656.17p 0 659.057p 0 659.058p 10000.0u 659.059p 0 659.447p 0 659.448p 10000.0u 659.449p 0 666.146p 0 666.147p 10000.0u 666.148p 0 678.914p 0 678.915p 10000.0u 678.916p 0 680.582p 0 680.583p 10000.0u 680.584p 0 698.933p 0 698.934p 10000.0u 698.935p 0 717.86p 0 717.861p 10000.0u 717.862p 0 721.46p 0 721.461p 10000.0u 721.462p 0 734.294p 0 734.295p 10000.0u 734.296p 0 740.642p 0 740.643p 10000.0u 740.644p 0 793.697p 0 793.698p 10000.0u 793.699p 0 797.159p 0 797.16p 10000.0u 797.161p 0 814.25p 0 814.251p 10000.0u 814.252p 0 824.894p 0 824.895p 10000.0u 824.896p 0 836.894p 0 836.895p 10000.0u 836.896p 0 842.579p 0 842.58p 10000.0u 842.581p 0 848.273p 0 848.274p 10000.0u 848.275p 0 850.898p 0 850.899p 10000.0u 850.9p 0 858.386p 0 858.387p 10000.0u 858.388p 0 868.925p 0 868.926p 10000.0u 868.927p 0 868.979p 0 868.98p 10000.0u 868.981p 0 877.718p 0 877.719p 10000.0u 877.72p 0 880.238p 0 880.239p 10000.0u 880.24p 0 881.993p 0 881.994p 10000.0u 881.995p 0 885.323p 0 885.324p 10000.0u 885.325p 0 913.373p 0 913.374p 10000.0u 913.375p 0 914.024p 0 914.025p 10000.0u 914.026p 0 923.768p 0 923.769p 10000.0u 923.77p 0 967.502p 0 967.503p 10000.0u 967.504p 0 978.221p 0 978.222p 10000.0u 978.223p 0 983.222p 0 983.223p 10000.0u 983.224p 0 992.108p 0 992.109p 10000.0u 992.11p 0 994.988p 0 994.989p 10000.0u 994.99p 0)
IIN86 0 87 pwl(0 0 12.269p 0 12.27p 10000.0u 12.271p 0 16.061p 0 16.062p 10000.0u 16.063p 0 20.336p 0 20.337p 10000.0u 20.338p 0 40.805p 0 40.806p 10000.0u 40.807p 0 50.807p 0 50.808p 10000.0u 50.809p 0 51.167p 0 51.168p 10000.0u 51.169p 0 51.635p 0 51.636p 10000.0u 51.637p 0 55.127p 0 55.128p 10000.0u 55.129p 0 65.252p 0 65.253p 10000.0u 65.254p 0 73.412p 0 73.413p 10000.0u 73.414p 0 78.257p 0 78.258p 10000.0u 78.259p 0 83.078p 0 83.079p 10000.0u 83.08p 0 89.666p 0 89.667p 10000.0u 89.668p 0 109.274p 0 109.275p 10000.0u 109.276p 0 121.181p 0 121.182p 10000.0u 121.183p 0 123.809p 0 123.81p 10000.0u 123.811p 0 124.472p 0 124.473p 10000.0u 124.474p 0 130.904p 0 130.905p 10000.0u 130.906p 0 160.664p 0 160.665p 10000.0u 160.666p 0 164.525p 0 164.526p 10000.0u 164.527p 0 175.907p 0 175.908p 10000.0u 175.909p 0 197.957p 0 197.958p 10000.0u 197.959p 0 205.172p 0 205.173p 10000.0u 205.174p 0 210.479p 0 210.48p 10000.0u 210.481p 0 211.742p 0 211.743p 10000.0u 211.744p 0 213.404p 0 213.405p 10000.0u 213.406p 0 247.805p 0 247.806p 10000.0u 247.807p 0 255.305p 0 255.306p 10000.0u 255.307p 0 278.561p 0 278.562p 10000.0u 278.563p 0 285.113p 0 285.114p 10000.0u 285.115p 0 285.752p 0 285.753p 10000.0u 285.754p 0 307.427p 0 307.428p 10000.0u 307.429p 0 313.415p 0 313.416p 10000.0u 313.417p 0 320.963p 0 320.964p 10000.0u 320.965p 0 333.659p 0 333.66p 10000.0u 333.661p 0 371.972p 0 371.973p 10000.0u 371.974p 0 372.572p 0 372.573p 10000.0u 372.574p 0 377.66p 0 377.661p 10000.0u 377.662p 0 383.648p 0 383.649p 10000.0u 383.65p 0 384.503p 0 384.504p 10000.0u 384.505p 0 387.806p 0 387.807p 10000.0u 387.808p 0 390.539p 0 390.54p 10000.0u 390.541p 0 416.576p 0 416.577p 10000.0u 416.578p 0 426.986p 0 426.987p 10000.0u 426.988p 0 442.121p 0 442.122p 10000.0u 442.123p 0 443.501p 0 443.502p 10000.0u 443.503p 0 445.409p 0 445.41p 10000.0u 445.411p 0 447.701p 0 447.702p 10000.0u 447.703p 0 449.627p 0 449.628p 10000.0u 449.629p 0 455.915p 0 455.916p 10000.0u 455.917p 0 462.773p 0 462.774p 10000.0u 462.775p 0 468.365p 0 468.366p 10000.0u 468.367p 0 486.068p 0 486.069p 10000.0u 486.07p 0 486.686p 0 486.687p 10000.0u 486.688p 0 517.43p 0 517.431p 10000.0u 517.432p 0 526.211p 0 526.212p 10000.0u 526.213p 0 531.098p 0 531.099p 10000.0u 531.1p 0 536.669p 0 536.67p 10000.0u 536.671p 0 537.677p 0 537.678p 10000.0u 537.679p 0 542.231p 0 542.232p 10000.0u 542.233p 0 545.678p 0 545.679p 10000.0u 545.68p 0 549.536p 0 549.537p 10000.0u 549.538p 0 552.566p 0 552.567p 10000.0u 552.568p 0 581.003p 0 581.004p 10000.0u 581.005p 0 587.888p 0 587.889p 10000.0u 587.89p 0 600.026p 0 600.027p 10000.0u 600.028p 0 602.804p 0 602.805p 10000.0u 602.806p 0 603.305p 0 603.306p 10000.0u 603.307p 0 609.836p 0 609.837p 10000.0u 609.838p 0 627.791p 0 627.792p 10000.0u 627.793p 0 638.105p 0 638.106p 10000.0u 638.107p 0 650.297p 0 650.298p 10000.0u 650.299p 0 659.669p 0 659.67p 10000.0u 659.671p 0 678.824p 0 678.825p 10000.0u 678.826p 0 696.305p 0 696.306p 10000.0u 696.307p 0 698.33p 0 698.331p 10000.0u 698.332p 0 707.165p 0 707.166p 10000.0u 707.167p 0 711.551p 0 711.552p 10000.0u 711.553p 0 713.09p 0 713.091p 10000.0u 713.092p 0 727.088p 0 727.089p 10000.0u 727.09p 0 732.278p 0 732.279p 10000.0u 732.28p 0 739.778p 0 739.779p 10000.0u 739.78p 0 742.316p 0 742.317p 10000.0u 742.318p 0 754.085p 0 754.086p 10000.0u 754.087p 0 755.915p 0 755.916p 10000.0u 755.917p 0 764.714p 0 764.715p 10000.0u 764.716p 0 765.977p 0 765.978p 10000.0u 765.979p 0 769.724p 0 769.725p 10000.0u 769.726p 0 770.747p 0 770.748p 10000.0u 770.749p 0 780.425p 0 780.426p 10000.0u 780.427p 0 791.75p 0 791.751p 10000.0u 791.752p 0 795.341p 0 795.342p 10000.0u 795.343p 0 798.284p 0 798.285p 10000.0u 798.286p 0 802.223p 0 802.224p 10000.0u 802.225p 0 821.87p 0 821.871p 10000.0u 821.872p 0 828.77p 0 828.771p 10000.0u 828.772p 0 829.016p 0 829.017p 10000.0u 829.018p 0 841.592p 0 841.593p 10000.0u 841.594p 0 856.259p 0 856.26p 10000.0u 856.261p 0 859.829p 0 859.83p 10000.0u 859.831p 0 863.912p 0 863.913p 10000.0u 863.914p 0 876.5p 0 876.501p 10000.0u 876.502p 0 916.013p 0 916.014p 10000.0u 916.015p 0 916.379p 0 916.38p 10000.0u 916.381p 0 946.61p 0 946.611p 10000.0u 946.612p 0 954.113p 0 954.114p 10000.0u 954.115p 0 957.632p 0 957.633p 10000.0u 957.634p 0 960.233p 0 960.234p 10000.0u 960.235p 0 974.702p 0 974.703p 10000.0u 974.704p 0)
IIN87 0 88 pwl(0 0 9.98p 0 9.981p 10000.0u 9.982p 0 22.28p 0 22.281p 10000.0u 22.282p 0 41.414p 0 41.415p 10000.0u 41.416p 0 54.14p 0 54.141p 10000.0u 54.142p 0 83.366p 0 83.367p 10000.0u 83.368p 0 91.073p 0 91.074p 10000.0u 91.075p 0 96.065p 0 96.066p 10000.0u 96.067p 0 97.553p 0 97.554p 10000.0u 97.555p 0 101.045p 0 101.046p 10000.0u 101.047p 0 103.838p 0 103.839p 10000.0u 103.84p 0 121.34p 0 121.341p 10000.0u 121.342p 0 126.395p 0 126.396p 10000.0u 126.397p 0 129.938p 0 129.939p 10000.0u 129.94p 0 135.902p 0 135.903p 10000.0u 135.904p 0 141.344p 0 141.345p 10000.0u 141.346p 0 142.469p 0 142.47p 10000.0u 142.471p 0 162.044p 0 162.045p 10000.0u 162.046p 0 162.623p 0 162.624p 10000.0u 162.625p 0 194.348p 0 194.349p 10000.0u 194.35p 0 206.324p 0 206.325p 10000.0u 206.326p 0 213.383p 0 213.384p 10000.0u 213.385p 0 216.785p 0 216.786p 10000.0u 216.787p 0 221.015p 0 221.016p 10000.0u 221.017p 0 222.953p 0 222.954p 10000.0u 222.955p 0 223.136p 0 223.137p 10000.0u 223.138p 0 223.658p 0 223.659p 10000.0u 223.66p 0 236.501p 0 236.502p 10000.0u 236.503p 0 240.473p 0 240.474p 10000.0u 240.475p 0 252.275p 0 252.276p 10000.0u 252.277p 0 259.046p 0 259.047p 10000.0u 259.048p 0 269.258p 0 269.259p 10000.0u 269.26p 0 276.242p 0 276.243p 10000.0u 276.244p 0 279.902p 0 279.903p 10000.0u 279.904p 0 281.399p 0 281.4p 10000.0u 281.401p 0 295.955p 0 295.956p 10000.0u 295.957p 0 299.657p 0 299.658p 10000.0u 299.659p 0 303.083p 0 303.084p 10000.0u 303.085p 0 333.17p 0 333.171p 10000.0u 333.172p 0 337.73p 0 337.731p 10000.0u 337.732p 0 348.443p 0 348.444p 10000.0u 348.445p 0 350.792p 0 350.793p 10000.0u 350.794p 0 353.333p 0 353.334p 10000.0u 353.335p 0 363.068p 0 363.069p 10000.0u 363.07p 0 367.031p 0 367.032p 10000.0u 367.033p 0 370.757p 0 370.758p 10000.0u 370.759p 0 372.206p 0 372.207p 10000.0u 372.208p 0 375.38p 0 375.381p 10000.0u 375.382p 0 385.616p 0 385.617p 10000.0u 385.618p 0 386.705p 0 386.706p 10000.0u 386.707p 0 395.009p 0 395.01p 10000.0u 395.011p 0 400.976p 0 400.977p 10000.0u 400.978p 0 402.356p 0 402.357p 10000.0u 402.358p 0 406.352p 0 406.353p 10000.0u 406.354p 0 424.865p 0 424.866p 10000.0u 424.867p 0 440.69p 0 440.691p 10000.0u 440.692p 0 441.542p 0 441.543p 10000.0u 441.544p 0 448.775p 0 448.776p 10000.0u 448.777p 0 449.549p 0 449.55p 10000.0u 449.551p 0 474.455p 0 474.456p 10000.0u 474.457p 0 502.472p 0 502.473p 10000.0u 502.474p 0 507.935p 0 507.936p 10000.0u 507.937p 0 529.829p 0 529.83p 10000.0u 529.831p 0 553.271p 0 553.272p 10000.0u 553.273p 0 641.075p 0 641.076p 10000.0u 641.077p 0 645.392p 0 645.393p 10000.0u 645.394p 0 654.623p 0 654.624p 10000.0u 654.625p 0 660.044p 0 660.045p 10000.0u 660.046p 0 675.485p 0 675.486p 10000.0u 675.487p 0 678.284p 0 678.285p 10000.0u 678.286p 0 681.56p 0 681.561p 10000.0u 681.562p 0 683.045p 0 683.046p 10000.0u 683.047p 0 683.789p 0 683.79p 10000.0u 683.791p 0 688.793p 0 688.794p 10000.0u 688.795p 0 709.364p 0 709.365p 10000.0u 709.366p 0 711.794p 0 711.795p 10000.0u 711.796p 0 712.793p 0 712.794p 10000.0u 712.795p 0 715.67p 0 715.671p 10000.0u 715.672p 0 717.701p 0 717.702p 10000.0u 717.703p 0 724.268p 0 724.269p 10000.0u 724.27p 0 725.231p 0 725.232p 10000.0u 725.233p 0 753.215p 0 753.216p 10000.0u 753.217p 0 762.776p 0 762.777p 10000.0u 762.778p 0 770.369p 0 770.37p 10000.0u 770.371p 0 783.89p 0 783.891p 10000.0u 783.892p 0 789.437p 0 789.438p 10000.0u 789.439p 0 790.964p 0 790.965p 10000.0u 790.966p 0 811.112p 0 811.113p 10000.0u 811.114p 0 829.238p 0 829.239p 10000.0u 829.24p 0 833.87p 0 833.871p 10000.0u 833.872p 0 857.501p 0 857.502p 10000.0u 857.503p 0 863.066p 0 863.067p 10000.0u 863.068p 0 898.916p 0 898.917p 10000.0u 898.918p 0 922.79p 0 922.791p 10000.0u 922.792p 0 926.132p 0 926.133p 10000.0u 926.134p 0 943.181p 0 943.182p 10000.0u 943.183p 0 945.503p 0 945.504p 10000.0u 945.505p 0 953.276p 0 953.277p 10000.0u 953.278p 0 986.108p 0 986.109p 10000.0u 986.11p 0 989.549p 0 989.55p 10000.0u 989.551p 0)
IIN88 0 89 pwl(0 0 9.566p 0 9.567p 10000.0u 9.568p 0 22.277p 0 22.278p 10000.0u 22.279p 0 32.348p 0 32.349p 10000.0u 32.35p 0 45.227p 0 45.228p 10000.0u 45.229p 0 50.741p 0 50.742p 10000.0u 50.743p 0 61.913p 0 61.914p 10000.0u 61.915p 0 63.32p 0 63.321p 10000.0u 63.322p 0 64.442p 0 64.443p 10000.0u 64.444p 0 66.584p 0 66.585p 10000.0u 66.586p 0 71.738p 0 71.739p 10000.0u 71.74p 0 77.915p 0 77.916p 10000.0u 77.917p 0 100.211p 0 100.212p 10000.0u 100.213p 0 103.436p 0 103.437p 10000.0u 103.438p 0 116.111p 0 116.112p 10000.0u 116.113p 0 116.627p 0 116.628p 10000.0u 116.629p 0 124.556p 0 124.557p 10000.0u 124.558p 0 131.945p 0 131.946p 10000.0u 131.947p 0 151.919p 0 151.92p 10000.0u 151.921p 0 158.462p 0 158.463p 10000.0u 158.464p 0 166.391p 0 166.392p 10000.0u 166.393p 0 173.387p 0 173.388p 10000.0u 173.389p 0 178.628p 0 178.629p 10000.0u 178.63p 0 187.922p 0 187.923p 10000.0u 187.924p 0 194.108p 0 194.109p 10000.0u 194.11p 0 195.86p 0 195.861p 10000.0u 195.862p 0 197.522p 0 197.523p 10000.0u 197.524p 0 214.382p 0 214.383p 10000.0u 214.384p 0 219.314p 0 219.315p 10000.0u 219.316p 0 230.897p 0 230.898p 10000.0u 230.899p 0 234.344p 0 234.345p 10000.0u 234.346p 0 247.202p 0 247.203p 10000.0u 247.204p 0 273.881p 0 273.882p 10000.0u 273.883p 0 281.936p 0 281.937p 10000.0u 281.938p 0 296.909p 0 296.91p 10000.0u 296.911p 0 305.159p 0 305.16p 10000.0u 305.161p 0 331.835p 0 331.836p 10000.0u 331.837p 0 343.133p 0 343.134p 10000.0u 343.135p 0 354.899p 0 354.9p 10000.0u 354.901p 0 355.133p 0 355.134p 10000.0u 355.135p 0 356.261p 0 356.262p 10000.0u 356.263p 0 371.483p 0 371.484p 10000.0u 371.485p 0 382.97p 0 382.971p 10000.0u 382.972p 0 387.131p 0 387.132p 10000.0u 387.133p 0 401.939p 0 401.94p 10000.0u 401.941p 0 409.241p 0 409.242p 10000.0u 409.243p 0 432.914p 0 432.915p 10000.0u 432.916p 0 433.145p 0 433.146p 10000.0u 433.147p 0 436.019p 0 436.02p 10000.0u 436.021p 0 440.081p 0 440.082p 10000.0u 440.083p 0 452.375p 0 452.376p 10000.0u 452.377p 0 471.968p 0 471.969p 10000.0u 471.97p 0 474.173p 0 474.174p 10000.0u 474.175p 0 482.357p 0 482.358p 10000.0u 482.359p 0 486.476p 0 486.477p 10000.0u 486.478p 0 512.192p 0 512.193p 10000.0u 512.194p 0 520.235p 0 520.236p 10000.0u 520.237p 0 540.137p 0 540.138p 10000.0u 540.139p 0 548.708p 0 548.709p 10000.0u 548.71p 0 570.374p 0 570.375p 10000.0u 570.376p 0 588.707p 0 588.708p 10000.0u 588.709p 0 592.697p 0 592.698p 10000.0u 592.699p 0 593.363p 0 593.364p 10000.0u 593.365p 0 593.612p 0 593.613p 10000.0u 593.614p 0 606.956p 0 606.957p 10000.0u 606.958p 0 614.651p 0 614.652p 10000.0u 614.653p 0 622.124p 0 622.125p 10000.0u 622.126p 0 625.754p 0 625.755p 10000.0u 625.756p 0 627.737p 0 627.738p 10000.0u 627.739p 0 640.772p 0 640.773p 10000.0u 640.774p 0 645.59p 0 645.591p 10000.0u 645.592p 0 658.34p 0 658.341p 10000.0u 658.342p 0 675.11p 0 675.111p 10000.0u 675.112p 0 676.721p 0 676.722p 10000.0u 676.723p 0 681.122p 0 681.123p 10000.0u 681.124p 0 685.664p 0 685.665p 10000.0u 685.666p 0 696.35p 0 696.351p 10000.0u 696.352p 0 697.865p 0 697.866p 10000.0u 697.867p 0 715.205p 0 715.206p 10000.0u 715.207p 0 723.431p 0 723.432p 10000.0u 723.433p 0 748.58p 0 748.581p 10000.0u 748.582p 0 792.383p 0 792.384p 10000.0u 792.385p 0 801.458p 0 801.459p 10000.0u 801.46p 0 806.453p 0 806.454p 10000.0u 806.455p 0 813.614p 0 813.615p 10000.0u 813.616p 0 833.723p 0 833.724p 10000.0u 833.725p 0 840.617p 0 840.618p 10000.0u 840.619p 0 849.647p 0 849.648p 10000.0u 849.649p 0 863.381p 0 863.382p 10000.0u 863.383p 0 878.816p 0 878.817p 10000.0u 878.818p 0 891.551p 0 891.552p 10000.0u 891.553p 0 910.403p 0 910.404p 10000.0u 910.405p 0 919.697p 0 919.698p 10000.0u 919.699p 0 920.102p 0 920.103p 10000.0u 920.104p 0 921.668p 0 921.669p 10000.0u 921.67p 0 956.864p 0 956.865p 10000.0u 956.866p 0 959.738p 0 959.739p 10000.0u 959.74p 0 967.469p 0 967.47p 10000.0u 967.471p 0 981.818p 0 981.819p 10000.0u 981.82p 0)
IIN89 0 90 pwl(0 0 9.311p 0 9.312p 10000.0u 9.313p 0 24.467p 0 24.468p 10000.0u 24.469p 0 24.803p 0 24.804p 10000.0u 24.805p 0 27.647p 0 27.648p 10000.0u 27.649p 0 44.597p 0 44.598p 10000.0u 44.599p 0 47.468p 0 47.469p 10000.0u 47.47p 0 48.65p 0 48.651p 10000.0u 48.652p 0 54.026p 0 54.027p 10000.0u 54.028p 0 55.562p 0 55.563p 10000.0u 55.564p 0 65.849p 0 65.85p 10000.0u 65.851p 0 69.398p 0 69.399p 10000.0u 69.4p 0 81.71p 0 81.711p 10000.0u 81.712p 0 86.627p 0 86.628p 10000.0u 86.629p 0 90.185p 0 90.186p 10000.0u 90.187p 0 94.127p 0 94.128p 10000.0u 94.129p 0 98.33p 0 98.331p 10000.0u 98.332p 0 107.741p 0 107.742p 10000.0u 107.743p 0 111.539p 0 111.54p 10000.0u 111.541p 0 128.633p 0 128.634p 10000.0u 128.635p 0 141.53p 0 141.531p 10000.0u 141.532p 0 143.024p 0 143.025p 10000.0u 143.026p 0 150.113p 0 150.114p 10000.0u 150.115p 0 150.845p 0 150.846p 10000.0u 150.847p 0 162.032p 0 162.033p 10000.0u 162.034p 0 178.865p 0 178.866p 10000.0u 178.867p 0 197.6p 0 197.601p 10000.0u 197.602p 0 206.549p 0 206.55p 10000.0u 206.551p 0 208.424p 0 208.425p 10000.0u 208.426p 0 217.751p 0 217.752p 10000.0u 217.753p 0 234.68p 0 234.681p 10000.0u 234.682p 0 235.136p 0 235.137p 10000.0u 235.138p 0 237.947p 0 237.948p 10000.0u 237.949p 0 271.745p 0 271.746p 10000.0u 271.747p 0 274.817p 0 274.818p 10000.0u 274.819p 0 289.571p 0 289.572p 10000.0u 289.573p 0 297.149p 0 297.15p 10000.0u 297.151p 0 298.298p 0 298.299p 10000.0u 298.3p 0 301.85p 0 301.851p 10000.0u 301.852p 0 310.751p 0 310.752p 10000.0u 310.753p 0 319.868p 0 319.869p 10000.0u 319.87p 0 337.643p 0 337.644p 10000.0u 337.645p 0 338.864p 0 338.865p 10000.0u 338.866p 0 342.344p 0 342.345p 10000.0u 342.346p 0 356.339p 0 356.34p 10000.0u 356.341p 0 384.938p 0 384.939p 10000.0u 384.94p 0 393.623p 0 393.624p 10000.0u 393.625p 0 396.512p 0 396.513p 10000.0u 396.514p 0 402.002p 0 402.003p 10000.0u 402.004p 0 403.16p 0 403.161p 10000.0u 403.162p 0 424.574p 0 424.575p 10000.0u 424.576p 0 451.838p 0 451.839p 10000.0u 451.84p 0 461.099p 0 461.1p 10000.0u 461.101p 0 475.883p 0 475.884p 10000.0u 475.885p 0 478.445p 0 478.446p 10000.0u 478.447p 0 478.934p 0 478.935p 10000.0u 478.936p 0 480.182p 0 480.183p 10000.0u 480.184p 0 489.332p 0 489.333p 10000.0u 489.334p 0 491.093p 0 491.094p 10000.0u 491.095p 0 494.405p 0 494.406p 10000.0u 494.407p 0 497.048p 0 497.049p 10000.0u 497.05p 0 499.262p 0 499.263p 10000.0u 499.264p 0 501.881p 0 501.882p 10000.0u 501.883p 0 509.72p 0 509.721p 10000.0u 509.722p 0 516.449p 0 516.45p 10000.0u 516.451p 0 530.435p 0 530.436p 10000.0u 530.437p 0 544.787p 0 544.788p 10000.0u 544.789p 0 552.386p 0 552.387p 10000.0u 552.388p 0 557.828p 0 557.829p 10000.0u 557.83p 0 573.794p 0 573.795p 10000.0u 573.796p 0 580.208p 0 580.209p 10000.0u 580.21p 0 585.701p 0 585.702p 10000.0u 585.703p 0 596.318p 0 596.319p 10000.0u 596.32p 0 603.944p 0 603.945p 10000.0u 603.946p 0 611.096p 0 611.097p 10000.0u 611.098p 0 615.821p 0 615.822p 10000.0u 615.823p 0 619.907p 0 619.908p 10000.0u 619.909p 0 650.246p 0 650.247p 10000.0u 650.248p 0 654.239p 0 654.24p 10000.0u 654.241p 0 663.608p 0 663.609p 10000.0u 663.61p 0 686.261p 0 686.262p 10000.0u 686.263p 0 696.821p 0 696.822p 10000.0u 696.823p 0 702.941p 0 702.942p 10000.0u 702.943p 0 707.549p 0 707.55p 10000.0u 707.551p 0 709.313p 0 709.314p 10000.0u 709.315p 0 714.779p 0 714.78p 10000.0u 714.781p 0 715.46p 0 715.461p 10000.0u 715.462p 0 723.971p 0 723.972p 10000.0u 723.973p 0 725.261p 0 725.262p 10000.0u 725.263p 0 785.774p 0 785.775p 10000.0u 785.776p 0 786.803p 0 786.804p 10000.0u 786.805p 0 788.129p 0 788.13p 10000.0u 788.131p 0 790.907p 0 790.908p 10000.0u 790.909p 0 797.63p 0 797.631p 10000.0u 797.632p 0 804.038p 0 804.039p 10000.0u 804.04p 0 821.318p 0 821.319p 10000.0u 821.32p 0 821.87p 0 821.871p 10000.0u 821.872p 0 830.216p 0 830.217p 10000.0u 830.218p 0 875.006p 0 875.007p 10000.0u 875.008p 0 876.308p 0 876.309p 10000.0u 876.31p 0 917.993p 0 917.994p 10000.0u 917.995p 0 925.445p 0 925.446p 10000.0u 925.447p 0 933.479p 0 933.48p 10000.0u 933.481p 0 937.931p 0 937.932p 10000.0u 937.933p 0 951.878p 0 951.879p 10000.0u 951.88p 0 953.852p 0 953.853p 10000.0u 953.854p 0 958.028p 0 958.029p 10000.0u 958.03p 0 960.977p 0 960.978p 10000.0u 960.979p 0 973.343p 0 973.344p 10000.0u 973.345p 0 981.596p 0 981.597p 10000.0u 981.598p 0 987.053p 0 987.054p 10000.0u 987.055p 0 991.37p 0 991.371p 10000.0u 991.372p 0 994.958p 0 994.959p 10000.0u 994.96p 0 997.013p 0 997.014p 10000.0u 997.015p 0)
IIN90 0 91 pwl(0 0 5.885p 0 5.886p 10000.0u 5.887p 0 13.859p 0 13.86p 10000.0u 13.861p 0 35.009p 0 35.01p 10000.0u 35.011p 0 39.83p 0 39.831p 10000.0u 39.832p 0 52.172p 0 52.173p 10000.0u 52.174p 0 52.832p 0 52.833p 10000.0u 52.834p 0 57.749p 0 57.75p 10000.0u 57.751p 0 60.485p 0 60.486p 10000.0u 60.487p 0 66.137p 0 66.138p 10000.0u 66.139p 0 91.466p 0 91.467p 10000.0u 91.468p 0 93.272p 0 93.273p 10000.0u 93.274p 0 100.784p 0 100.785p 10000.0u 100.786p 0 106.121p 0 106.122p 10000.0u 106.123p 0 160.352p 0 160.353p 10000.0u 160.354p 0 175.706p 0 175.707p 10000.0u 175.708p 0 186.299p 0 186.3p 10000.0u 186.301p 0 187.046p 0 187.047p 10000.0u 187.048p 0 240.395p 0 240.396p 10000.0u 240.397p 0 243.437p 0 243.438p 10000.0u 243.439p 0 265.763p 0 265.764p 10000.0u 265.765p 0 268.688p 0 268.689p 10000.0u 268.69p 0 302.234p 0 302.235p 10000.0u 302.236p 0 305.165p 0 305.166p 10000.0u 305.167p 0 320.231p 0 320.232p 10000.0u 320.233p 0 324.989p 0 324.99p 10000.0u 324.991p 0 333.842p 0 333.843p 10000.0u 333.844p 0 335.534p 0 335.535p 10000.0u 335.536p 0 341.726p 0 341.727p 10000.0u 341.728p 0 355.556p 0 355.557p 10000.0u 355.558p 0 380.093p 0 380.094p 10000.0u 380.095p 0 391.364p 0 391.365p 10000.0u 391.366p 0 401.213p 0 401.214p 10000.0u 401.215p 0 405.743p 0 405.744p 10000.0u 405.745p 0 435.656p 0 435.657p 10000.0u 435.658p 0 439.34p 0 439.341p 10000.0u 439.342p 0 439.619p 0 439.62p 10000.0u 439.621p 0 443.822p 0 443.823p 10000.0u 443.824p 0 463.682p 0 463.683p 10000.0u 463.684p 0 466.814p 0 466.815p 10000.0u 466.816p 0 479.378p 0 479.379p 10000.0u 479.38p 0 505.604p 0 505.605p 10000.0u 505.606p 0 512.474p 0 512.475p 10000.0u 512.476p 0 524.303p 0 524.304p 10000.0u 524.305p 0 526.172p 0 526.173p 10000.0u 526.174p 0 528.197p 0 528.198p 10000.0u 528.199p 0 541.421p 0 541.422p 10000.0u 541.423p 0 545.321p 0 545.322p 10000.0u 545.323p 0 568.124p 0 568.125p 10000.0u 568.126p 0 574.961p 0 574.962p 10000.0u 574.963p 0 587.942p 0 587.943p 10000.0u 587.944p 0 591.926p 0 591.927p 10000.0u 591.928p 0 604.148p 0 604.149p 10000.0u 604.15p 0 625.334p 0 625.335p 10000.0u 625.336p 0 648.638p 0 648.639p 10000.0u 648.64p 0 649.937p 0 649.938p 10000.0u 649.939p 0 652.934p 0 652.935p 10000.0u 652.936p 0 683.264p 0 683.265p 10000.0u 683.266p 0 704.054p 0 704.055p 10000.0u 704.056p 0 717.341p 0 717.342p 10000.0u 717.343p 0 743.327p 0 743.328p 10000.0u 743.329p 0 746.063p 0 746.064p 10000.0u 746.065p 0 751.151p 0 751.152p 10000.0u 751.153p 0 767.174p 0 767.175p 10000.0u 767.176p 0 770.078p 0 770.079p 10000.0u 770.08p 0 774.092p 0 774.093p 10000.0u 774.094p 0 800.63p 0 800.631p 10000.0u 800.632p 0 807.14p 0 807.141p 10000.0u 807.142p 0 817.133p 0 817.134p 10000.0u 817.135p 0 844.286p 0 844.287p 10000.0u 844.288p 0 856.775p 0 856.776p 10000.0u 856.777p 0 885.659p 0 885.66p 10000.0u 885.661p 0 892.592p 0 892.593p 10000.0u 892.594p 0 911.195p 0 911.196p 10000.0u 911.197p 0 911.876p 0 911.877p 10000.0u 911.878p 0 922.781p 0 922.782p 10000.0u 922.783p 0 926.711p 0 926.712p 10000.0u 926.713p 0 943.157p 0 943.158p 10000.0u 943.159p 0 946.013p 0 946.014p 10000.0u 946.015p 0 954.683p 0 954.684p 10000.0u 954.685p 0 964.541p 0 964.542p 10000.0u 964.543p 0 966.557p 0 966.558p 10000.0u 966.559p 0 969.737p 0 969.738p 10000.0u 969.739p 0 975.935p 0 975.936p 10000.0u 975.937p 0 982.949p 0 982.95p 10000.0u 982.951p 0 983.621p 0 983.622p 10000.0u 983.623p 0 991.937p 0 991.938p 10000.0u 991.939p 0 992.438p 0 992.439p 10000.0u 992.44p 0 999.377p 0 999.378p 10000.0u 999.379p 0 999.854p 0 999.855p 10000.0u 999.856p 0)
IIN91 0 92 pwl(0 0 7.697p 0 7.698p 10000.0u 7.699p 0 10.982p 0 10.983p 10000.0u 10.984p 0 12.926p 0 12.927p 10000.0u 12.928p 0 23.402p 0 23.403p 10000.0u 23.404p 0 24.407p 0 24.408p 10000.0u 24.409p 0 30.671p 0 30.672p 10000.0u 30.673p 0 36.287p 0 36.288p 10000.0u 36.289p 0 37.382p 0 37.383p 10000.0u 37.384p 0 41.147p 0 41.148p 10000.0u 41.149p 0 53.567p 0 53.568p 10000.0u 53.569p 0 54.623p 0 54.624p 10000.0u 54.625p 0 58.028p 0 58.029p 10000.0u 58.03p 0 71.435p 0 71.436p 10000.0u 71.437p 0 75.671p 0 75.672p 10000.0u 75.673p 0 79.544p 0 79.545p 10000.0u 79.546p 0 81.152p 0 81.153p 10000.0u 81.154p 0 93.206p 0 93.207p 10000.0u 93.208p 0 130.982p 0 130.983p 10000.0u 130.984p 0 133.349p 0 133.35p 10000.0u 133.351p 0 140.987p 0 140.988p 10000.0u 140.989p 0 147.857p 0 147.858p 10000.0u 147.859p 0 171.92p 0 171.921p 10000.0u 171.922p 0 173.039p 0 173.04p 10000.0u 173.041p 0 176.018p 0 176.019p 10000.0u 176.02p 0 190.412p 0 190.413p 10000.0u 190.414p 0 225.806p 0 225.807p 10000.0u 225.808p 0 230.525p 0 230.526p 10000.0u 230.527p 0 243.134p 0 243.135p 10000.0u 243.136p 0 249.203p 0 249.204p 10000.0u 249.205p 0 252.818p 0 252.819p 10000.0u 252.82p 0 254.432p 0 254.433p 10000.0u 254.434p 0 259.976p 0 259.977p 10000.0u 259.978p 0 270.344p 0 270.345p 10000.0u 270.346p 0 285.878p 0 285.879p 10000.0u 285.88p 0 305.405p 0 305.406p 10000.0u 305.407p 0 309.728p 0 309.729p 10000.0u 309.73p 0 325.238p 0 325.239p 10000.0u 325.24p 0 340.241p 0 340.242p 10000.0u 340.243p 0 346.259p 0 346.26p 10000.0u 346.261p 0 355.178p 0 355.179p 10000.0u 355.18p 0 366.224p 0 366.225p 10000.0u 366.226p 0 367.484p 0 367.485p 10000.0u 367.486p 0 373.748p 0 373.749p 10000.0u 373.75p 0 382.88p 0 382.881p 10000.0u 382.882p 0 386.216p 0 386.217p 10000.0u 386.218p 0 389.129p 0 389.13p 10000.0u 389.131p 0 389.186p 0 389.187p 10000.0u 389.188p 0 391.148p 0 391.149p 10000.0u 391.15p 0 400.01p 0 400.011p 10000.0u 400.012p 0 416.606p 0 416.607p 10000.0u 416.608p 0 417.908p 0 417.909p 10000.0u 417.91p 0 419.657p 0 419.658p 10000.0u 419.659p 0 425.495p 0 425.496p 10000.0u 425.497p 0 444.935p 0 444.936p 10000.0u 444.937p 0 448.319p 0 448.32p 10000.0u 448.321p 0 474.29p 0 474.291p 10000.0u 474.292p 0 503.783p 0 503.784p 10000.0u 503.785p 0 506.552p 0 506.553p 10000.0u 506.554p 0 514.604p 0 514.605p 10000.0u 514.606p 0 522.395p 0 522.396p 10000.0u 522.397p 0 533.333p 0 533.334p 10000.0u 533.335p 0 547.76p 0 547.761p 10000.0u 547.762p 0 554.519p 0 554.52p 10000.0u 554.521p 0 573.929p 0 573.93p 10000.0u 573.931p 0 606.725p 0 606.726p 10000.0u 606.727p 0 614.747p 0 614.748p 10000.0u 614.749p 0 624.932p 0 624.933p 10000.0u 624.934p 0 627.83p 0 627.831p 10000.0u 627.832p 0 652.895p 0 652.896p 10000.0u 652.897p 0 655.217p 0 655.218p 10000.0u 655.219p 0 659.714p 0 659.715p 10000.0u 659.716p 0 669.257p 0 669.258p 10000.0u 669.259p 0 681.932p 0 681.933p 10000.0u 681.934p 0 694.808p 0 694.809p 10000.0u 694.81p 0 698.027p 0 698.028p 10000.0u 698.029p 0 702.71p 0 702.711p 10000.0u 702.712p 0 712.433p 0 712.434p 10000.0u 712.435p 0 713.099p 0 713.1p 10000.0u 713.101p 0 727.658p 0 727.659p 10000.0u 727.66p 0 730.835p 0 730.836p 10000.0u 730.837p 0 732.782p 0 732.783p 10000.0u 732.784p 0 733.247p 0 733.248p 10000.0u 733.249p 0 745.04p 0 745.041p 10000.0u 745.042p 0 754.421p 0 754.422p 10000.0u 754.423p 0 768.875p 0 768.876p 10000.0u 768.877p 0 775.958p 0 775.959p 10000.0u 775.96p 0 779.396p 0 779.397p 10000.0u 779.398p 0 801.185p 0 801.186p 10000.0u 801.187p 0 805.037p 0 805.038p 10000.0u 805.039p 0 810.986p 0 810.987p 10000.0u 810.988p 0 823.43p 0 823.431p 10000.0u 823.432p 0 825.929p 0 825.93p 10000.0u 825.931p 0 832.883p 0 832.884p 10000.0u 832.885p 0 866.735p 0 866.736p 10000.0u 866.737p 0 867.833p 0 867.834p 10000.0u 867.835p 0 868.97p 0 868.971p 10000.0u 868.972p 0 888.023p 0 888.024p 10000.0u 888.025p 0 894.872p 0 894.873p 10000.0u 894.874p 0 898.691p 0 898.692p 10000.0u 898.693p 0 926.978p 0 926.979p 10000.0u 926.98p 0 944.711p 0 944.712p 10000.0u 944.713p 0 945.137p 0 945.138p 10000.0u 945.139p 0 983.339p 0 983.34p 10000.0u 983.341p 0 985.049p 0 985.05p 10000.0u 985.051p 0 985.418p 0 985.419p 10000.0u 985.42p 0 998.444p 0 998.445p 10000.0u 998.446p 0)
IIN92 0 93 pwl(0 0 5.75p 0 5.751p 10000.0u 5.752p 0 25.547p 0 25.548p 10000.0u 25.549p 0 27.548p 0 27.549p 10000.0u 27.55p 0 47.387p 0 47.388p 10000.0u 47.389p 0 52.346p 0 52.347p 10000.0u 52.348p 0 54.797p 0 54.798p 10000.0u 54.799p 0 64.742p 0 64.743p 10000.0u 64.744p 0 73.544p 0 73.545p 10000.0u 73.546p 0 83.237p 0 83.238p 10000.0u 83.239p 0 89.219p 0 89.22p 10000.0u 89.221p 0 100.175p 0 100.176p 10000.0u 100.177p 0 100.733p 0 100.734p 10000.0u 100.735p 0 105.791p 0 105.792p 10000.0u 105.793p 0 116.195p 0 116.196p 10000.0u 116.197p 0 118.247p 0 118.248p 10000.0u 118.249p 0 126.158p 0 126.159p 10000.0u 126.16p 0 128.906p 0 128.907p 10000.0u 128.908p 0 139.058p 0 139.059p 10000.0u 139.06p 0 144.359p 0 144.36p 10000.0u 144.361p 0 158.933p 0 158.934p 10000.0u 158.935p 0 164.852p 0 164.853p 10000.0u 164.854p 0 176.234p 0 176.235p 10000.0u 176.236p 0 202.451p 0 202.452p 10000.0u 202.453p 0 213.545p 0 213.546p 10000.0u 213.547p 0 220.001p 0 220.002p 10000.0u 220.003p 0 228.155p 0 228.156p 10000.0u 228.157p 0 230.21p 0 230.211p 10000.0u 230.212p 0 243.866p 0 243.867p 10000.0u 243.868p 0 244.229p 0 244.23p 10000.0u 244.231p 0 246.269p 0 246.27p 10000.0u 246.271p 0 254.003p 0 254.004p 10000.0u 254.005p 0 271.22p 0 271.221p 10000.0u 271.222p 0 272.618p 0 272.619p 10000.0u 272.62p 0 284.072p 0 284.073p 10000.0u 284.074p 0 300.938p 0 300.939p 10000.0u 300.94p 0 321.989p 0 321.99p 10000.0u 321.991p 0 327.284p 0 327.285p 10000.0u 327.286p 0 334.805p 0 334.806p 10000.0u 334.807p 0 337.772p 0 337.773p 10000.0u 337.774p 0 339.728p 0 339.729p 10000.0u 339.73p 0 341.897p 0 341.898p 10000.0u 341.899p 0 348.869p 0 348.87p 10000.0u 348.871p 0 372.548p 0 372.549p 10000.0u 372.55p 0 384.617p 0 384.618p 10000.0u 384.619p 0 385.874p 0 385.875p 10000.0u 385.876p 0 411.332p 0 411.333p 10000.0u 411.334p 0 430.28p 0 430.281p 10000.0u 430.282p 0 436.652p 0 436.653p 10000.0u 436.654p 0 457.931p 0 457.932p 10000.0u 457.933p 0 461.777p 0 461.778p 10000.0u 461.779p 0 467.144p 0 467.145p 10000.0u 467.146p 0 469.139p 0 469.14p 10000.0u 469.141p 0 494.483p 0 494.484p 10000.0u 494.485p 0 501.35p 0 501.351p 10000.0u 501.352p 0 508.517p 0 508.518p 10000.0u 508.519p 0 522.233p 0 522.234p 10000.0u 522.235p 0 527.054p 0 527.055p 10000.0u 527.056p 0 528.254p 0 528.255p 10000.0u 528.256p 0 533.39p 0 533.391p 10000.0u 533.392p 0 534.176p 0 534.177p 10000.0u 534.178p 0 534.629p 0 534.63p 10000.0u 534.631p 0 548.555p 0 548.556p 10000.0u 548.557p 0 550.004p 0 550.005p 10000.0u 550.006p 0 551.078p 0 551.079p 10000.0u 551.08p 0 553.481p 0 553.482p 10000.0u 553.483p 0 554.591p 0 554.592p 10000.0u 554.593p 0 575.126p 0 575.127p 10000.0u 575.128p 0 578.852p 0 578.853p 10000.0u 578.854p 0 586.565p 0 586.566p 10000.0u 586.567p 0 598.403p 0 598.404p 10000.0u 598.405p 0 603.167p 0 603.168p 10000.0u 603.169p 0 607.433p 0 607.434p 10000.0u 607.435p 0 619.409p 0 619.41p 10000.0u 619.411p 0 647.348p 0 647.349p 10000.0u 647.35p 0 653.036p 0 653.037p 10000.0u 653.038p 0 659.648p 0 659.649p 10000.0u 659.65p 0 666.989p 0 666.99p 10000.0u 666.991p 0 689.84p 0 689.841p 10000.0u 689.842p 0 707.663p 0 707.664p 10000.0u 707.665p 0 731.258p 0 731.259p 10000.0u 731.26p 0 743.369p 0 743.37p 10000.0u 743.371p 0 746.207p 0 746.208p 10000.0u 746.209p 0 748.211p 0 748.212p 10000.0u 748.213p 0 754.103p 0 754.104p 10000.0u 754.105p 0 760.805p 0 760.806p 10000.0u 760.807p 0 768.344p 0 768.345p 10000.0u 768.346p 0 778.067p 0 778.068p 10000.0u 778.069p 0 782.915p 0 782.916p 10000.0u 782.917p 0 793.424p 0 793.425p 10000.0u 793.426p 0 810.179p 0 810.18p 10000.0u 810.181p 0 823.133p 0 823.134p 10000.0u 823.135p 0 830.636p 0 830.637p 10000.0u 830.638p 0 840.164p 0 840.165p 10000.0u 840.166p 0 851.321p 0 851.322p 10000.0u 851.323p 0 859.361p 0 859.362p 10000.0u 859.363p 0 862.373p 0 862.374p 10000.0u 862.375p 0 873.2p 0 873.201p 10000.0u 873.202p 0 882.29p 0 882.291p 10000.0u 882.292p 0 885.557p 0 885.558p 10000.0u 885.559p 0 894.272p 0 894.273p 10000.0u 894.274p 0 895.274p 0 895.275p 10000.0u 895.276p 0 907.457p 0 907.458p 10000.0u 907.459p 0 908.459p 0 908.46p 10000.0u 908.461p 0 915.803p 0 915.804p 10000.0u 915.805p 0 920.144p 0 920.145p 10000.0u 920.146p 0 926.339p 0 926.34p 10000.0u 926.341p 0 952.331p 0 952.332p 10000.0u 952.333p 0 966.821p 0 966.822p 10000.0u 966.823p 0 969.008p 0 969.009p 10000.0u 969.01p 0 973.151p 0 973.152p 10000.0u 973.153p 0 981.743p 0 981.744p 10000.0u 981.745p 0 982.313p 0 982.314p 10000.0u 982.315p 0 982.883p 0 982.884p 10000.0u 982.885p 0 994.832p 0 994.833p 10000.0u 994.834p 0)
IIN93 0 94 pwl(0 0 1.967p 0 1.968p 10000.0u 1.969p 0 2.813p 0 2.814p 10000.0u 2.815p 0 11.957p 0 11.958p 10000.0u 11.959p 0 13.337p 0 13.338p 10000.0u 13.339p 0 23.789p 0 23.79p 10000.0u 23.791p 0 26.276p 0 26.277p 10000.0u 26.278p 0 26.537p 0 26.538p 10000.0u 26.539p 0 33.065p 0 33.066p 10000.0u 33.067p 0 36.308p 0 36.309p 10000.0u 36.31p 0 39.809p 0 39.81p 10000.0u 39.811p 0 42.074p 0 42.075p 10000.0u 42.076p 0 45.515p 0 45.516p 10000.0u 45.517p 0 61.523p 0 61.524p 10000.0u 61.525p 0 70.676p 0 70.677p 10000.0u 70.678p 0 77.0p 0 77.001p 10000.0u 77.002p 0 85.4p 0 85.401p 10000.0u 85.402p 0 98.267p 0 98.268p 10000.0u 98.269p 0 108.917p 0 108.918p 10000.0u 108.919p 0 109.601p 0 109.602p 10000.0u 109.603p 0 111.917p 0 111.918p 10000.0u 111.919p 0 116.975p 0 116.976p 10000.0u 116.977p 0 126.539p 0 126.54p 10000.0u 126.541p 0 149.819p 0 149.82p 10000.0u 149.821p 0 154.94p 0 154.941p 10000.0u 154.942p 0 165.293p 0 165.294p 10000.0u 165.295p 0 192.575p 0 192.576p 10000.0u 192.577p 0 192.794p 0 192.795p 10000.0u 192.796p 0 193.067p 0 193.068p 10000.0u 193.069p 0 203.036p 0 203.037p 10000.0u 203.038p 0 203.414p 0 203.415p 10000.0u 203.416p 0 206.762p 0 206.763p 10000.0u 206.764p 0 232.076p 0 232.077p 10000.0u 232.078p 0 236.996p 0 236.997p 10000.0u 236.998p 0 238.037p 0 238.038p 10000.0u 238.039p 0 246.428p 0 246.429p 10000.0u 246.43p 0 262.223p 0 262.224p 10000.0u 262.225p 0 271.808p 0 271.809p 10000.0u 271.81p 0 290.003p 0 290.004p 10000.0u 290.005p 0 298.307p 0 298.308p 10000.0u 298.309p 0 307.955p 0 307.956p 10000.0u 307.957p 0 316.559p 0 316.56p 10000.0u 316.561p 0 325.286p 0 325.287p 10000.0u 325.288p 0 333.323p 0 333.324p 10000.0u 333.325p 0 354.677p 0 354.678p 10000.0u 354.679p 0 368.792p 0 368.793p 10000.0u 368.794p 0 370.169p 0 370.17p 10000.0u 370.171p 0 377.054p 0 377.055p 10000.0u 377.056p 0 404.492p 0 404.493p 10000.0u 404.494p 0 441.86p 0 441.861p 10000.0u 441.862p 0 442.964p 0 442.965p 10000.0u 442.966p 0 451.091p 0 451.092p 10000.0u 451.093p 0 466.211p 0 466.212p 10000.0u 466.213p 0 468.017p 0 468.018p 10000.0u 468.019p 0 469.295p 0 469.296p 10000.0u 469.297p 0 470.279p 0 470.28p 10000.0u 470.281p 0 485.714p 0 485.715p 10000.0u 485.716p 0 486.221p 0 486.222p 10000.0u 486.223p 0 511.685p 0 511.686p 10000.0u 511.687p 0 513.926p 0 513.927p 10000.0u 513.928p 0 526.466p 0 526.467p 10000.0u 526.468p 0 532.295p 0 532.296p 10000.0u 532.297p 0 539.222p 0 539.223p 10000.0u 539.224p 0 545.765p 0 545.766p 10000.0u 545.767p 0 549.284p 0 549.285p 10000.0u 549.286p 0 555.59p 0 555.591p 10000.0u 555.592p 0 564.683p 0 564.684p 10000.0u 564.685p 0 569.063p 0 569.064p 10000.0u 569.065p 0 585.83p 0 585.831p 10000.0u 585.832p 0 614.138p 0 614.139p 10000.0u 614.14p 0 621.434p 0 621.435p 10000.0u 621.436p 0 626.72p 0 626.721p 10000.0u 626.722p 0 644.168p 0 644.169p 10000.0u 644.17p 0 650.135p 0 650.136p 10000.0u 650.137p 0 655.775p 0 655.776p 10000.0u 655.777p 0 656.444p 0 656.445p 10000.0u 656.446p 0 672.371p 0 672.372p 10000.0u 672.373p 0 676.994p 0 676.995p 10000.0u 676.996p 0 679.838p 0 679.839p 10000.0u 679.84p 0 680.948p 0 680.949p 10000.0u 680.95p 0 685.463p 0 685.464p 10000.0u 685.465p 0 695.237p 0 695.238p 10000.0u 695.239p 0 702.212p 0 702.213p 10000.0u 702.214p 0 709.904p 0 709.905p 10000.0u 709.906p 0 714.911p 0 714.912p 10000.0u 714.913p 0 722.711p 0 722.712p 10000.0u 722.713p 0 725.792p 0 725.793p 10000.0u 725.794p 0 738.734p 0 738.735p 10000.0u 738.736p 0 744.329p 0 744.33p 10000.0u 744.331p 0 748.85p 0 748.851p 10000.0u 748.852p 0 769.808p 0 769.809p 10000.0u 769.81p 0 785.507p 0 785.508p 10000.0u 785.509p 0 795.293p 0 795.294p 10000.0u 795.295p 0 832.706p 0 832.707p 10000.0u 832.708p 0 835.181p 0 835.182p 10000.0u 835.183p 0 842.69p 0 842.691p 10000.0u 842.692p 0 854.444p 0 854.445p 10000.0u 854.446p 0 854.789p 0 854.79p 10000.0u 854.791p 0 876.77p 0 876.771p 10000.0u 876.772p 0 883.754p 0 883.755p 10000.0u 883.756p 0 893.354p 0 893.355p 10000.0u 893.356p 0 893.405p 0 893.406p 10000.0u 893.407p 0 899.816p 0 899.817p 10000.0u 899.818p 0 914.99p 0 914.991p 10000.0u 914.992p 0 919.295p 0 919.296p 10000.0u 919.297p 0 926.432p 0 926.433p 10000.0u 926.434p 0 948.278p 0 948.279p 10000.0u 948.28p 0 951.524p 0 951.525p 10000.0u 951.526p 0 957.722p 0 957.723p 10000.0u 957.724p 0 959.867p 0 959.868p 10000.0u 959.869p 0 962.519p 0 962.52p 10000.0u 962.521p 0 972.386p 0 972.387p 10000.0u 972.388p 0 973.832p 0 973.833p 10000.0u 973.834p 0 978.419p 0 978.42p 10000.0u 978.421p 0 981.971p 0 981.972p 10000.0u 981.973p 0 984.755p 0 984.756p 10000.0u 984.757p 0)
IIN94 0 95 pwl(0 0 7.925p 0 7.926p 10000.0u 7.927p 0 18.266p 0 18.267p 10000.0u 18.268p 0 31.982p 0 31.983p 10000.0u 31.984p 0 42.455p 0 42.456p 10000.0u 42.457p 0 46.514p 0 46.515p 10000.0u 46.516p 0 54.215p 0 54.216p 10000.0u 54.217p 0 58.829p 0 58.83p 10000.0u 58.831p 0 67.967p 0 67.968p 10000.0u 67.969p 0 68.6p 0 68.601p 10000.0u 68.602p 0 77.69p 0 77.691p 10000.0u 77.692p 0 80.63p 0 80.631p 10000.0u 80.632p 0 103.124p 0 103.125p 10000.0u 103.126p 0 104.75p 0 104.751p 10000.0u 104.752p 0 107.735p 0 107.736p 10000.0u 107.737p 0 119.807p 0 119.808p 10000.0u 119.809p 0 133.541p 0 133.542p 10000.0u 133.543p 0 140.759p 0 140.76p 10000.0u 140.761p 0 141.344p 0 141.345p 10000.0u 141.346p 0 146.942p 0 146.943p 10000.0u 146.944p 0 148.352p 0 148.353p 10000.0u 148.354p 0 150.866p 0 150.867p 10000.0u 150.868p 0 154.718p 0 154.719p 10000.0u 154.72p 0 185.141p 0 185.142p 10000.0u 185.143p 0 187.292p 0 187.293p 10000.0u 187.294p 0 191.285p 0 191.286p 10000.0u 191.287p 0 198.782p 0 198.783p 10000.0u 198.784p 0 202.592p 0 202.593p 10000.0u 202.594p 0 235.592p 0 235.593p 10000.0u 235.594p 0 242.525p 0 242.526p 10000.0u 242.527p 0 243.206p 0 243.207p 10000.0u 243.208p 0 256.334p 0 256.335p 10000.0u 256.336p 0 258.722p 0 258.723p 10000.0u 258.724p 0 260.633p 0 260.634p 10000.0u 260.635p 0 262.307p 0 262.308p 10000.0u 262.309p 0 265.379p 0 265.38p 10000.0u 265.381p 0 283.01p 0 283.011p 10000.0u 283.012p 0 295.175p 0 295.176p 10000.0u 295.177p 0 299.153p 0 299.154p 10000.0u 299.155p 0 299.309p 0 299.31p 10000.0u 299.311p 0 299.735p 0 299.736p 10000.0u 299.737p 0 305.459p 0 305.46p 10000.0u 305.461p 0 312.659p 0 312.66p 10000.0u 312.661p 0 314.42p 0 314.421p 10000.0u 314.422p 0 319.811p 0 319.812p 10000.0u 319.813p 0 335.276p 0 335.277p 10000.0u 335.278p 0 346.523p 0 346.524p 10000.0u 346.525p 0 351.578p 0 351.579p 10000.0u 351.58p 0 359.471p 0 359.472p 10000.0u 359.473p 0 378.401p 0 378.402p 10000.0u 378.403p 0 426.629p 0 426.63p 10000.0u 426.631p 0 429.353p 0 429.354p 10000.0u 429.355p 0 435.212p 0 435.213p 10000.0u 435.214p 0 447.233p 0 447.234p 10000.0u 447.235p 0 454.127p 0 454.128p 10000.0u 454.129p 0 459.233p 0 459.234p 10000.0u 459.235p 0 464.675p 0 464.676p 10000.0u 464.677p 0 466.955p 0 466.956p 10000.0u 466.957p 0 470.825p 0 470.826p 10000.0u 470.827p 0 471.617p 0 471.618p 10000.0u 471.619p 0 471.845p 0 471.846p 10000.0u 471.847p 0 474.116p 0 474.117p 10000.0u 474.118p 0 486.665p 0 486.666p 10000.0u 486.667p 0 488.771p 0 488.772p 10000.0u 488.773p 0 495.017p 0 495.018p 10000.0u 495.019p 0 498.878p 0 498.879p 10000.0u 498.88p 0 504.569p 0 504.57p 10000.0u 504.571p 0 515.447p 0 515.448p 10000.0u 515.449p 0 518.321p 0 518.322p 10000.0u 518.323p 0 523.292p 0 523.293p 10000.0u 523.294p 0 533.369p 0 533.37p 10000.0u 533.371p 0 541.475p 0 541.476p 10000.0u 541.477p 0 550.247p 0 550.248p 10000.0u 550.249p 0 553.904p 0 553.905p 10000.0u 553.906p 0 553.916p 0 553.917p 10000.0u 553.918p 0 559.391p 0 559.392p 10000.0u 559.393p 0 561.788p 0 561.789p 10000.0u 561.79p 0 571.145p 0 571.146p 10000.0u 571.147p 0 588.878p 0 588.879p 10000.0u 588.88p 0 593.297p 0 593.298p 10000.0u 593.299p 0 605.372p 0 605.373p 10000.0u 605.374p 0 621.095p 0 621.096p 10000.0u 621.097p 0 622.529p 0 622.53p 10000.0u 622.531p 0 636.338p 0 636.339p 10000.0u 636.34p 0 642.056p 0 642.057p 10000.0u 642.058p 0 656.738p 0 656.739p 10000.0u 656.74p 0 665.831p 0 665.832p 10000.0u 665.833p 0 669.836p 0 669.837p 10000.0u 669.838p 0 686.291p 0 686.292p 10000.0u 686.293p 0 697.091p 0 697.092p 10000.0u 697.093p 0 700.427p 0 700.428p 10000.0u 700.429p 0 705.437p 0 705.438p 10000.0u 705.439p 0 747.554p 0 747.555p 10000.0u 747.556p 0 748.19p 0 748.191p 10000.0u 748.192p 0 755.759p 0 755.76p 10000.0u 755.761p 0 783.095p 0 783.096p 10000.0u 783.097p 0 785.147p 0 785.148p 10000.0u 785.149p 0 804.743p 0 804.744p 10000.0u 804.745p 0 808.352p 0 808.353p 10000.0u 808.354p 0 813.566p 0 813.567p 10000.0u 813.568p 0 816.131p 0 816.132p 10000.0u 816.133p 0 816.785p 0 816.786p 10000.0u 816.787p 0 816.917p 0 816.918p 10000.0u 816.919p 0 821.777p 0 821.778p 10000.0u 821.779p 0 822.686p 0 822.687p 10000.0u 822.688p 0 824.126p 0 824.127p 10000.0u 824.128p 0 824.966p 0 824.967p 10000.0u 824.968p 0 838.535p 0 838.536p 10000.0u 838.537p 0 843.605p 0 843.606p 10000.0u 843.607p 0 845.717p 0 845.718p 10000.0u 845.719p 0 852.605p 0 852.606p 10000.0u 852.607p 0 869.459p 0 869.46p 10000.0u 869.461p 0 883.331p 0 883.332p 10000.0u 883.333p 0 886.52p 0 886.521p 10000.0u 886.522p 0 905.942p 0 905.943p 10000.0u 905.944p 0 913.406p 0 913.407p 10000.0u 913.408p 0 933.419p 0 933.42p 10000.0u 933.421p 0 946.451p 0 946.452p 10000.0u 946.453p 0 946.979p 0 946.98p 10000.0u 946.981p 0 949.589p 0 949.59p 10000.0u 949.591p 0 963.749p 0 963.75p 10000.0u 963.751p 0 976.52p 0 976.521p 10000.0u 976.522p 0 995.732p 0 995.733p 10000.0u 995.734p 0 997.958p 0 997.959p 10000.0u 997.96p 0 999.407p 0 999.408p 10000.0u 999.409p 0)
IIN95 0 96 pwl(0 0 27.047p 0 27.048p 10000.0u 27.049p 0 36.488p 0 36.489p 10000.0u 36.49p 0 67.106p 0 67.107p 10000.0u 67.108p 0 67.193p 0 67.194p 10000.0u 67.195p 0 106.604p 0 106.605p 10000.0u 106.606p 0 113.414p 0 113.415p 10000.0u 113.416p 0 116.099p 0 116.1p 10000.0u 116.101p 0 120.434p 0 120.435p 10000.0u 120.436p 0 134.201p 0 134.202p 10000.0u 134.203p 0 149.243p 0 149.244p 10000.0u 149.245p 0 155.966p 0 155.967p 10000.0u 155.968p 0 163.199p 0 163.2p 10000.0u 163.201p 0 163.841p 0 163.842p 10000.0u 163.843p 0 165.023p 0 165.024p 10000.0u 165.025p 0 165.53p 0 165.531p 10000.0u 165.532p 0 174.443p 0 174.444p 10000.0u 174.445p 0 187.4p 0 187.401p 10000.0u 187.402p 0 195.602p 0 195.603p 10000.0u 195.604p 0 201.953p 0 201.954p 10000.0u 201.955p 0 230.279p 0 230.28p 10000.0u 230.281p 0 243.311p 0 243.312p 10000.0u 243.313p 0 298.55p 0 298.551p 10000.0u 298.552p 0 301.367p 0 301.368p 10000.0u 301.369p 0 334.196p 0 334.197p 10000.0u 334.198p 0 338.654p 0 338.655p 10000.0u 338.656p 0 348.095p 0 348.096p 10000.0u 348.097p 0 388.832p 0 388.833p 10000.0u 388.834p 0 399.932p 0 399.933p 10000.0u 399.934p 0 400.61p 0 400.611p 10000.0u 400.612p 0 412.394p 0 412.395p 10000.0u 412.396p 0 412.667p 0 412.668p 10000.0u 412.669p 0 425.042p 0 425.043p 10000.0u 425.044p 0 440.645p 0 440.646p 10000.0u 440.647p 0 442.949p 0 442.95p 10000.0u 442.951p 0 445.187p 0 445.188p 10000.0u 445.189p 0 469.901p 0 469.902p 10000.0u 469.903p 0 482.729p 0 482.73p 10000.0u 482.731p 0 487.694p 0 487.695p 10000.0u 487.696p 0 494.183p 0 494.184p 10000.0u 494.185p 0 495.317p 0 495.318p 10000.0u 495.319p 0 505.403p 0 505.404p 10000.0u 505.405p 0 506.351p 0 506.352p 10000.0u 506.353p 0 529.562p 0 529.563p 10000.0u 529.564p 0 549.779p 0 549.78p 10000.0u 549.781p 0 556.229p 0 556.23p 10000.0u 556.231p 0 566.612p 0 566.613p 10000.0u 566.614p 0 587.69p 0 587.691p 10000.0u 587.692p 0 593.063p 0 593.064p 10000.0u 593.065p 0 602.6p 0 602.601p 10000.0u 602.602p 0 610.61p 0 610.611p 10000.0u 610.612p 0 617.255p 0 617.256p 10000.0u 617.257p 0 622.562p 0 622.563p 10000.0u 622.564p 0 623.276p 0 623.277p 10000.0u 623.278p 0 642.554p 0 642.555p 10000.0u 642.556p 0 649.721p 0 649.722p 10000.0u 649.723p 0 653.0p 0 653.001p 10000.0u 653.002p 0 661.169p 0 661.17p 10000.0u 661.171p 0 662.39p 0 662.391p 10000.0u 662.392p 0 679.106p 0 679.107p 10000.0u 679.108p 0 683.771p 0 683.772p 10000.0u 683.773p 0 714.776p 0 714.777p 10000.0u 714.778p 0 721.082p 0 721.083p 10000.0u 721.084p 0 740.618p 0 740.619p 10000.0u 740.62p 0 756.707p 0 756.708p 10000.0u 756.709p 0 758.441p 0 758.442p 10000.0u 758.443p 0 767.873p 0 767.874p 10000.0u 767.875p 0 796.553p 0 796.554p 10000.0u 796.555p 0 797.774p 0 797.775p 10000.0u 797.776p 0 808.7p 0 808.701p 10000.0u 808.702p 0 824.612p 0 824.613p 10000.0u 824.614p 0 825.902p 0 825.903p 10000.0u 825.904p 0 840.857p 0 840.858p 10000.0u 840.859p 0 876.386p 0 876.387p 10000.0u 876.388p 0 877.904p 0 877.905p 10000.0u 877.906p 0 885.512p 0 885.513p 10000.0u 885.514p 0 890.129p 0 890.13p 10000.0u 890.131p 0 899.72p 0 899.721p 10000.0u 899.722p 0 900.359p 0 900.36p 10000.0u 900.361p 0 903.275p 0 903.276p 10000.0u 903.277p 0 909.056p 0 909.057p 10000.0u 909.058p 0 917.924p 0 917.925p 10000.0u 917.926p 0 933.806p 0 933.807p 10000.0u 933.808p 0 953.465p 0 953.466p 10000.0u 953.467p 0 955.391p 0 955.392p 10000.0u 955.393p 0 980.48p 0 980.481p 10000.0u 980.482p 0 981.566p 0 981.567p 10000.0u 981.568p 0 985.511p 0 985.512p 10000.0u 985.513p 0 988.217p 0 988.218p 10000.0u 988.219p 0)
IIN96 0 97 pwl(0 0 1.163p 0 1.164p 10000.0u 1.165p 0 14.753p 0 14.754p 10000.0u 14.755p 0 16.22p 0 16.221p 10000.0u 16.222p 0 26.03p 0 26.031p 10000.0u 26.032p 0 30.614p 0 30.615p 10000.0u 30.616p 0 35.597p 0 35.598p 10000.0u 35.599p 0 37.103p 0 37.104p 10000.0u 37.105p 0 43.196p 0 43.197p 10000.0u 43.198p 0 44.015p 0 44.016p 10000.0u 44.017p 0 48.434p 0 48.435p 10000.0u 48.436p 0 61.619p 0 61.62p 10000.0u 61.621p 0 67.811p 0 67.812p 10000.0u 67.813p 0 73.586p 0 73.587p 10000.0u 73.588p 0 80.039p 0 80.04p 10000.0u 80.041p 0 84.866p 0 84.867p 10000.0u 84.868p 0 88.013p 0 88.014p 10000.0u 88.015p 0 104.186p 0 104.187p 10000.0u 104.188p 0 104.297p 0 104.298p 10000.0u 104.299p 0 111.731p 0 111.732p 10000.0u 111.733p 0 151.631p 0 151.632p 10000.0u 151.633p 0 154.028p 0 154.029p 10000.0u 154.03p 0 156.383p 0 156.384p 10000.0u 156.385p 0 170.384p 0 170.385p 10000.0u 170.386p 0 186.917p 0 186.918p 10000.0u 186.919p 0 232.727p 0 232.728p 10000.0u 232.729p 0 233.966p 0 233.967p 10000.0u 233.968p 0 242.441p 0 242.442p 10000.0u 242.443p 0 249.89p 0 249.891p 10000.0u 249.892p 0 259.916p 0 259.917p 10000.0u 259.918p 0 276.806p 0 276.807p 10000.0u 276.808p 0 277.946p 0 277.947p 10000.0u 277.948p 0 279.122p 0 279.123p 10000.0u 279.124p 0 311.12p 0 311.121p 10000.0u 311.122p 0 312.545p 0 312.546p 10000.0u 312.547p 0 329.417p 0 329.418p 10000.0u 329.419p 0 333.71p 0 333.711p 10000.0u 333.712p 0 334.841p 0 334.842p 10000.0u 334.843p 0 344.432p 0 344.433p 10000.0u 344.434p 0 347.618p 0 347.619p 10000.0u 347.62p 0 350.012p 0 350.013p 10000.0u 350.014p 0 372.092p 0 372.093p 10000.0u 372.094p 0 395.282p 0 395.283p 10000.0u 395.284p 0 399.809p 0 399.81p 10000.0u 399.811p 0 410.783p 0 410.784p 10000.0u 410.785p 0 411.788p 0 411.789p 10000.0u 411.79p 0 425.006p 0 425.007p 10000.0u 425.008p 0 426.506p 0 426.507p 10000.0u 426.508p 0 426.512p 0 426.513p 10000.0u 426.514p 0 434.429p 0 434.43p 10000.0u 434.431p 0 437.948p 0 437.949p 10000.0u 437.95p 0 438.137p 0 438.138p 10000.0u 438.139p 0 451.484p 0 451.485p 10000.0u 451.486p 0 463.997p 0 463.998p 10000.0u 463.999p 0 481.715p 0 481.716p 10000.0u 481.717p 0 503.318p 0 503.319p 10000.0u 503.32p 0 520.997p 0 520.998p 10000.0u 520.999p 0 524.486p 0 524.487p 10000.0u 524.488p 0 538.934p 0 538.935p 10000.0u 538.936p 0 568.817p 0 568.818p 10000.0u 568.819p 0 577.316p 0 577.317p 10000.0u 577.318p 0 582.905p 0 582.906p 10000.0u 582.907p 0 584.135p 0 584.136p 10000.0u 584.137p 0 585.677p 0 585.678p 10000.0u 585.679p 0 593.663p 0 593.664p 10000.0u 593.665p 0 598.367p 0 598.368p 10000.0u 598.369p 0 600.281p 0 600.282p 10000.0u 600.283p 0 612.017p 0 612.018p 10000.0u 612.019p 0 623.195p 0 623.196p 10000.0u 623.197p 0 624.311p 0 624.312p 10000.0u 624.313p 0 631.523p 0 631.524p 10000.0u 631.525p 0 637.679p 0 637.68p 10000.0u 637.681p 0 646.166p 0 646.167p 10000.0u 646.168p 0 682.592p 0 682.593p 10000.0u 682.594p 0 683.153p 0 683.154p 10000.0u 683.155p 0 694.712p 0 694.713p 10000.0u 694.714p 0 695.885p 0 695.886p 10000.0u 695.887p 0 713.153p 0 713.154p 10000.0u 713.155p 0 713.528p 0 713.529p 10000.0u 713.53p 0 720.236p 0 720.237p 10000.0u 720.238p 0 723.158p 0 723.159p 10000.0u 723.16p 0 742.982p 0 742.983p 10000.0u 742.984p 0 752.879p 0 752.88p 10000.0u 752.881p 0 756.584p 0 756.585p 10000.0u 756.586p 0 769.532p 0 769.533p 10000.0u 769.534p 0 774.761p 0 774.762p 10000.0u 774.763p 0 782.669p 0 782.67p 10000.0u 782.671p 0 798.608p 0 798.609p 10000.0u 798.61p 0 799.331p 0 799.332p 10000.0u 799.333p 0 810.554p 0 810.555p 10000.0u 810.556p 0 821.21p 0 821.211p 10000.0u 821.212p 0 837.209p 0 837.21p 10000.0u 837.211p 0 847.784p 0 847.785p 10000.0u 847.786p 0 872.09p 0 872.091p 10000.0u 872.092p 0 910.922p 0 910.923p 10000.0u 910.924p 0 937.037p 0 937.038p 10000.0u 937.039p 0 995.687p 0 995.688p 10000.0u 995.689p 0 999.62p 0 999.621p 10000.0u 999.622p 0)
IIN97 0 98 pwl(0 0 28.898p 0 28.899p 10000.0u 28.9p 0 37.835p 0 37.836p 10000.0u 37.837p 0 50.201p 0 50.202p 10000.0u 50.203p 0 50.237p 0 50.238p 10000.0u 50.239p 0 60.056p 0 60.057p 10000.0u 60.058p 0 62.975p 0 62.976p 10000.0u 62.977p 0 64.148p 0 64.149p 10000.0u 64.15p 0 73.874p 0 73.875p 10000.0u 73.876p 0 86.855p 0 86.856p 10000.0u 86.857p 0 93.245p 0 93.246p 10000.0u 93.247p 0 101.393p 0 101.394p 10000.0u 101.395p 0 117.701p 0 117.702p 10000.0u 117.703p 0 119.654p 0 119.655p 10000.0u 119.656p 0 122.099p 0 122.1p 10000.0u 122.101p 0 134.105p 0 134.106p 10000.0u 134.107p 0 140.756p 0 140.757p 10000.0u 140.758p 0 140.909p 0 140.91p 10000.0u 140.911p 0 154.997p 0 154.998p 10000.0u 154.999p 0 160.43p 0 160.431p 10000.0u 160.432p 0 169.361p 0 169.362p 10000.0u 169.363p 0 188.816p 0 188.817p 10000.0u 188.818p 0 210.221p 0 210.222p 10000.0u 210.223p 0 213.893p 0 213.894p 10000.0u 213.895p 0 250.577p 0 250.578p 10000.0u 250.579p 0 254.618p 0 254.619p 10000.0u 254.62p 0 261.458p 0 261.459p 10000.0u 261.46p 0 261.89p 0 261.891p 10000.0u 261.892p 0 280.193p 0 280.194p 10000.0u 280.195p 0 287.039p 0 287.04p 10000.0u 287.041p 0 288.395p 0 288.396p 10000.0u 288.397p 0 290.81p 0 290.811p 10000.0u 290.812p 0 300.992p 0 300.993p 10000.0u 300.994p 0 305.192p 0 305.193p 10000.0u 305.194p 0 355.169p 0 355.17p 10000.0u 355.171p 0 366.566p 0 366.567p 10000.0u 366.568p 0 366.863p 0 366.864p 10000.0u 366.865p 0 372.524p 0 372.525p 10000.0u 372.526p 0 374.603p 0 374.604p 10000.0u 374.605p 0 403.349p 0 403.35p 10000.0u 403.351p 0 404.651p 0 404.652p 10000.0u 404.653p 0 406.637p 0 406.638p 10000.0u 406.639p 0 409.643p 0 409.644p 10000.0u 409.645p 0 429.17p 0 429.171p 10000.0u 429.172p 0 434.474p 0 434.475p 10000.0u 434.476p 0 440.822p 0 440.823p 10000.0u 440.824p 0 445.688p 0 445.689p 10000.0u 445.69p 0 460.577p 0 460.578p 10000.0u 460.579p 0 465.923p 0 465.924p 10000.0u 465.925p 0 480.392p 0 480.393p 10000.0u 480.394p 0 480.551p 0 480.552p 10000.0u 480.553p 0 487.283p 0 487.284p 10000.0u 487.285p 0 488.996p 0 488.997p 10000.0u 488.998p 0 495.968p 0 495.969p 10000.0u 495.97p 0 505.091p 0 505.092p 10000.0u 505.093p 0 510.506p 0 510.507p 10000.0u 510.508p 0 511.877p 0 511.878p 10000.0u 511.879p 0 517.511p 0 517.512p 10000.0u 517.513p 0 531.857p 0 531.858p 10000.0u 531.859p 0 532.346p 0 532.347p 10000.0u 532.348p 0 548.126p 0 548.127p 10000.0u 548.128p 0 549.077p 0 549.078p 10000.0u 549.079p 0 550.82p 0 550.821p 10000.0u 550.822p 0 568.091p 0 568.092p 10000.0u 568.093p 0 591.644p 0 591.645p 10000.0u 591.646p 0 592.385p 0 592.386p 10000.0u 592.387p 0 618.917p 0 618.918p 10000.0u 618.919p 0 625.652p 0 625.653p 10000.0u 625.654p 0 645.245p 0 645.246p 10000.0u 645.247p 0 660.635p 0 660.636p 10000.0u 660.637p 0 672.074p 0 672.075p 10000.0u 672.076p 0 678.878p 0 678.879p 10000.0u 678.88p 0 681.233p 0 681.234p 10000.0u 681.235p 0 681.713p 0 681.714p 10000.0u 681.715p 0 685.571p 0 685.572p 10000.0u 685.573p 0 695.219p 0 695.22p 10000.0u 695.221p 0 729.827p 0 729.828p 10000.0u 729.829p 0 738.941p 0 738.942p 10000.0u 738.943p 0 740.303p 0 740.304p 10000.0u 740.305p 0 747.17p 0 747.171p 10000.0u 747.172p 0 751.154p 0 751.155p 10000.0u 751.156p 0 755.897p 0 755.898p 10000.0u 755.899p 0 770.348p 0 770.349p 10000.0u 770.35p 0 778.943p 0 778.944p 10000.0u 778.945p 0 779.729p 0 779.73p 10000.0u 779.731p 0 779.927p 0 779.928p 10000.0u 779.929p 0 781.247p 0 781.248p 10000.0u 781.249p 0 852.893p 0 852.894p 10000.0u 852.895p 0 853.685p 0 853.686p 10000.0u 853.687p 0 867.536p 0 867.537p 10000.0u 867.538p 0 885.524p 0 885.525p 10000.0u 885.526p 0 887.285p 0 887.286p 10000.0u 887.287p 0 888.239p 0 888.24p 10000.0u 888.241p 0 902.039p 0 902.04p 10000.0u 902.041p 0 904.112p 0 904.113p 10000.0u 904.114p 0 917.078p 0 917.079p 10000.0u 917.08p 0 926.732p 0 926.733p 10000.0u 926.734p 0 944.3p 0 944.301p 10000.0u 944.302p 0 969.107p 0 969.108p 10000.0u 969.109p 0 977.543p 0 977.544p 10000.0u 977.545p 0 978.662p 0 978.663p 10000.0u 978.664p 0)
IIN98 0 99 pwl(0 0 5.051p 0 5.052p 10000.0u 5.053p 0 8.831p 0 8.832p 10000.0u 8.833p 0 35.261p 0 35.262p 10000.0u 35.263p 0 39.662p 0 39.663p 10000.0u 39.664p 0 45.845p 0 45.846p 10000.0u 45.847p 0 48.143p 0 48.144p 10000.0u 48.145p 0 59.237p 0 59.238p 10000.0u 59.239p 0 68.405p 0 68.406p 10000.0u 68.407p 0 93.968p 0 93.969p 10000.0u 93.97p 0 104.039p 0 104.04p 10000.0u 104.041p 0 136.976p 0 136.977p 10000.0u 136.978p 0 141.416p 0 141.417p 10000.0u 141.418p 0 145.097p 0 145.098p 10000.0u 145.099p 0 149.042p 0 149.043p 10000.0u 149.044p 0 175.103p 0 175.104p 10000.0u 175.105p 0 192.527p 0 192.528p 10000.0u 192.529p 0 196.724p 0 196.725p 10000.0u 196.726p 0 208.556p 0 208.557p 10000.0u 208.558p 0 214.379p 0 214.38p 10000.0u 214.381p 0 234.764p 0 234.765p 10000.0u 234.766p 0 236.543p 0 236.544p 10000.0u 236.545p 0 242.837p 0 242.838p 10000.0u 242.839p 0 254.654p 0 254.655p 10000.0u 254.656p 0 261.233p 0 261.234p 10000.0u 261.235p 0 267.434p 0 267.435p 10000.0u 267.436p 0 314.042p 0 314.043p 10000.0u 314.044p 0 315.929p 0 315.93p 10000.0u 315.931p 0 321.395p 0 321.396p 10000.0u 321.397p 0 323.606p 0 323.607p 10000.0u 323.608p 0 328.493p 0 328.494p 10000.0u 328.495p 0 331.403p 0 331.404p 10000.0u 331.405p 0 345.797p 0 345.798p 10000.0u 345.799p 0 349.94p 0 349.941p 10000.0u 349.942p 0 353.297p 0 353.298p 10000.0u 353.299p 0 359.993p 0 359.994p 10000.0u 359.995p 0 361.037p 0 361.038p 10000.0u 361.039p 0 361.061p 0 361.062p 10000.0u 361.063p 0 378.92p 0 378.921p 10000.0u 378.922p 0 389.474p 0 389.475p 10000.0u 389.476p 0 395.318p 0 395.319p 10000.0u 395.32p 0 398.042p 0 398.043p 10000.0u 398.044p 0 412.229p 0 412.23p 10000.0u 412.231p 0 413.828p 0 413.829p 10000.0u 413.83p 0 423.716p 0 423.717p 10000.0u 423.718p 0 434.528p 0 434.529p 10000.0u 434.53p 0 439.988p 0 439.989p 10000.0u 439.99p 0 446.996p 0 446.997p 10000.0u 446.998p 0 453.782p 0 453.783p 10000.0u 453.784p 0 468.647p 0 468.648p 10000.0u 468.649p 0 471.353p 0 471.354p 10000.0u 471.355p 0 474.974p 0 474.975p 10000.0u 474.976p 0 507.599p 0 507.6p 10000.0u 507.601p 0 517.589p 0 517.59p 10000.0u 517.591p 0 521.996p 0 521.997p 10000.0u 521.998p 0 534.479p 0 534.48p 10000.0u 534.481p 0 535.262p 0 535.263p 10000.0u 535.264p 0 543.044p 0 543.045p 10000.0u 543.046p 0 546.104p 0 546.105p 10000.0u 546.106p 0 550.436p 0 550.437p 10000.0u 550.438p 0 554.78p 0 554.781p 10000.0u 554.782p 0 568.034p 0 568.035p 10000.0u 568.036p 0 593.678p 0 593.679p 10000.0u 593.68p 0 594.05p 0 594.051p 10000.0u 594.052p 0 598.202p 0 598.203p 10000.0u 598.204p 0 613.601p 0 613.602p 10000.0u 613.603p 0 618.443p 0 618.444p 10000.0u 618.445p 0 618.476p 0 618.477p 10000.0u 618.478p 0 620.729p 0 620.73p 10000.0u 620.731p 0 664.892p 0 664.893p 10000.0u 664.894p 0 671.207p 0 671.208p 10000.0u 671.209p 0 676.064p 0 676.065p 10000.0u 676.066p 0 677.405p 0 677.406p 10000.0u 677.407p 0 702.293p 0 702.294p 10000.0u 702.295p 0 712.973p 0 712.974p 10000.0u 712.975p 0 763.61p 0 763.611p 10000.0u 763.612p 0 765.959p 0 765.96p 10000.0u 765.961p 0 771.323p 0 771.324p 10000.0u 771.325p 0 784.505p 0 784.506p 10000.0u 784.507p 0 789.794p 0 789.795p 10000.0u 789.796p 0 815.48p 0 815.481p 10000.0u 815.482p 0 817.559p 0 817.56p 10000.0u 817.561p 0 825.938p 0 825.939p 10000.0u 825.94p 0 834.629p 0 834.63p 10000.0u 834.631p 0 838.397p 0 838.398p 10000.0u 838.399p 0 848.837p 0 848.838p 10000.0u 848.839p 0 863.453p 0 863.454p 10000.0u 863.455p 0 874.313p 0 874.314p 10000.0u 874.315p 0 885.038p 0 885.039p 10000.0u 885.04p 0 890.735p 0 890.736p 10000.0u 890.737p 0 890.771p 0 890.772p 10000.0u 890.773p 0 901.223p 0 901.224p 10000.0u 901.225p 0 907.625p 0 907.626p 10000.0u 907.627p 0 910.652p 0 910.653p 10000.0u 910.654p 0 914.327p 0 914.328p 10000.0u 914.329p 0 916.571p 0 916.572p 10000.0u 916.573p 0 923.165p 0 923.166p 10000.0u 923.167p 0 934.991p 0 934.992p 10000.0u 934.993p 0 937.148p 0 937.149p 10000.0u 937.15p 0 939.653p 0 939.654p 10000.0u 939.655p 0 967.49p 0 967.491p 10000.0u 967.492p 0 968.99p 0 968.991p 10000.0u 968.992p 0 983.402p 0 983.403p 10000.0u 983.404p 0 993.89p 0 993.891p 10000.0u 993.892p 0)
IIN99 0 100 pwl(0 0 0.374p 0 0.375p 10000.0u 0.376p 0 16.736p 0 16.737p 10000.0u 16.738p 0 44.093p 0 44.094p 10000.0u 44.095p 0 54.203p 0 54.204p 10000.0u 54.205p 0 65.636p 0 65.637p 10000.0u 65.638p 0 70.277p 0 70.278p 10000.0u 70.279p 0 71.846p 0 71.847p 10000.0u 71.848p 0 78.632p 0 78.633p 10000.0u 78.634p 0 81.44p 0 81.441p 10000.0u 81.442p 0 85.172p 0 85.173p 10000.0u 85.174p 0 105.254p 0 105.255p 10000.0u 105.256p 0 110.084p 0 110.085p 10000.0u 110.086p 0 110.636p 0 110.637p 10000.0u 110.638p 0 125.813p 0 125.814p 10000.0u 125.815p 0 134.699p 0 134.7p 10000.0u 134.701p 0 148.856p 0 148.857p 10000.0u 148.858p 0 153.197p 0 153.198p 10000.0u 153.199p 0 156.941p 0 156.942p 10000.0u 156.943p 0 166.262p 0 166.263p 10000.0u 166.264p 0 173.93p 0 173.931p 10000.0u 173.932p 0 187.115p 0 187.116p 10000.0u 187.117p 0 188.648p 0 188.649p 10000.0u 188.65p 0 189.548p 0 189.549p 10000.0u 189.55p 0 229.676p 0 229.677p 10000.0u 229.678p 0 232.544p 0 232.545p 10000.0u 232.546p 0 235.235p 0 235.236p 10000.0u 235.237p 0 237.119p 0 237.12p 10000.0u 237.121p 0 246.428p 0 246.429p 10000.0u 246.43p 0 255.461p 0 255.462p 10000.0u 255.463p 0 278.231p 0 278.232p 10000.0u 278.233p 0 294.287p 0 294.288p 10000.0u 294.289p 0 299.375p 0 299.376p 10000.0u 299.377p 0 300.923p 0 300.924p 10000.0u 300.925p 0 304.691p 0 304.692p 10000.0u 304.693p 0 318.806p 0 318.807p 10000.0u 318.808p 0 356.645p 0 356.646p 10000.0u 356.647p 0 370.52p 0 370.521p 10000.0u 370.522p 0 399.677p 0 399.678p 10000.0u 399.679p 0 404.738p 0 404.739p 10000.0u 404.74p 0 407.501p 0 407.502p 10000.0u 407.503p 0 413.195p 0 413.196p 10000.0u 413.197p 0 429.188p 0 429.189p 10000.0u 429.19p 0 447.665p 0 447.666p 10000.0u 447.667p 0 450.872p 0 450.873p 10000.0u 450.874p 0 464.264p 0 464.265p 10000.0u 464.266p 0 469.22p 0 469.221p 10000.0u 469.222p 0 474.497p 0 474.498p 10000.0u 474.499p 0 494.579p 0 494.58p 10000.0u 494.581p 0 502.244p 0 502.245p 10000.0u 502.246p 0 515.291p 0 515.292p 10000.0u 515.293p 0 534.431p 0 534.432p 10000.0u 534.433p 0 543.779p 0 543.78p 10000.0u 543.781p 0 554.375p 0 554.376p 10000.0u 554.377p 0 578.936p 0 578.937p 10000.0u 578.938p 0 585.563p 0 585.564p 10000.0u 585.565p 0 592.859p 0 592.86p 10000.0u 592.861p 0 613.463p 0 613.464p 10000.0u 613.465p 0 614.237p 0 614.238p 10000.0u 614.239p 0 637.019p 0 637.02p 10000.0u 637.021p 0 641.096p 0 641.097p 10000.0u 641.098p 0 678.152p 0 678.153p 10000.0u 678.154p 0 679.739p 0 679.74p 10000.0u 679.741p 0 682.502p 0 682.503p 10000.0u 682.504p 0 691.526p 0 691.527p 10000.0u 691.528p 0 693.023p 0 693.024p 10000.0u 693.025p 0 695.489p 0 695.49p 10000.0u 695.491p 0 721.742p 0 721.743p 10000.0u 721.744p 0 728.093p 0 728.094p 10000.0u 728.095p 0 734.228p 0 734.229p 10000.0u 734.23p 0 749.453p 0 749.454p 10000.0u 749.455p 0 761.945p 0 761.946p 10000.0u 761.947p 0 778.76p 0 778.761p 10000.0u 778.762p 0 784.436p 0 784.437p 10000.0u 784.438p 0 795.722p 0 795.723p 10000.0u 795.724p 0 799.382p 0 799.383p 10000.0u 799.384p 0 803.351p 0 803.352p 10000.0u 803.353p 0 808.802p 0 808.803p 10000.0u 808.804p 0 809.522p 0 809.523p 10000.0u 809.524p 0 813.872p 0 813.873p 10000.0u 813.874p 0 823.697p 0 823.698p 10000.0u 823.699p 0 839.009p 0 839.01p 10000.0u 839.011p 0 843.788p 0 843.789p 10000.0u 843.79p 0 847.466p 0 847.467p 10000.0u 847.468p 0 862.142p 0 862.143p 10000.0u 862.144p 0 875.564p 0 875.565p 10000.0u 875.566p 0 884.495p 0 884.496p 10000.0u 884.497p 0 888.338p 0 888.339p 10000.0u 888.34p 0 919.664p 0 919.665p 10000.0u 919.666p 0 936.668p 0 936.669p 10000.0u 936.67p 0 948.644p 0 948.645p 10000.0u 948.646p 0 949.124p 0 949.125p 10000.0u 949.126p 0 950.594p 0 950.595p 10000.0u 950.596p 0 952.19p 0 952.191p 10000.0u 952.192p 0 980.489p 0 980.49p 10000.0u 980.491p 0 983.774p 0 983.775p 10000.0u 983.776p 0)

X0 exc-neuron 0 1 58 88 56 53 86 62 72 14 20 85 
X1 exc-neuron 0 2 53 76 51 83 32 90 63 81 87 96 
X2 exc-neuron 0 3 66 38 73 36 95 82 90 10 4 85 
X3 exc-neuron 0 4 35 3 71 91 80 28 87 2 56 45 
X4 exc-neuron 0 5 78 29 66 43 25 61 48 71 3 86 
X5 exc-neuron 0 6 85 38 24 62 78 33 36 98 69 68 
X6 exc-neuron 0 7 11 65 63 34 70 69 53 89 36 79 
X7 exc-neuron 0 8 62 72 23 85 13 51 15 37 54 26 
X8 exc-neuron 0 9 98 50 29 32 46 96 57 21 89 39 
X9 exc-neuron 0 10 49 92 21 14 38 84 51 8 6 48 
X10 exc-neuron 0 11 44 93 55 74 43 10 1 59 45 72 
X11 exc-neuron 0 12 58 31 61 89 40 37 23 70 99 57 
X12 exc-neuron 0 13 55 41 9 48 35 59 78 16 47 2 
X13 exc-neuron 0 14 5 36 45 37 16 80 3 15 26 54 
X14 exc-neuron 0 15 54 18 98 64 31 77 10 37 75 7 
X15 exc-neuron 0 16 66 23 70 64 82 41 49 96 56 90 
X16 exc-neuron 0 17 87 44 7 50 93 94 38 10 65 16 
X17 exc-neuron 0 18 37 88 32 14 27 5 57 21 56 15 
X18 exc-neuron 0 19 65 46 94 16 43 57 62 84 96 12 
X19 exc-neuron 0 20 82 63 92 5 85 91 2 83 29 43 
X20 exc-neuron 0 21 9 32 68 94 58 35 70 62 41 6 
X21 exc-neuron 0 22 98 95 82 85 13 75 46 88 54 76 
X22 exc-neuron 0 23 68 43 30 92 79 3 18 32 6 95 
X23 exc-neuron 0 24 86 2 94 69 5 47 64 70 16 44 
X24 exc-neuron 0 25 32 46 7 88 79 66 65 75 59 74 
X25 exc-neuron 0 26 12 17 19 84 91 59 33 13 66 2 
X26 exc-neuron 0 27 39 54 11 12 67 92 31 43 81 3 
X27 exc-neuron 0 28 39 12 40 34 96 25 84 92 23 86 
X28 exc-neuron 0 29 84 49 45 63 55 36 25 67 74 89 
X29 exc-neuron 0 30 73 47 88 37 34 85 25 9 13 29 
X30 exc-neuron 0 31 15 89 94 30 32 92 4 7 67 83 
X31 exc-neuron 0 32 72 15 74 28 65 9 12 94 51 6 
X32 exc-neuron 0 33 55 61 60 100 7 41 93 81 30 34 
X33 exc-neuron 0 34 65 28 85 18 13 76 17 38 59 81 
X34 exc-neuron 0 35 6 83 59 73 45 62 79 49 38 50 
X35 exc-neuron 0 36 12 11 47 41 24 60 62 37 52 4 
X36 exc-neuron 0 37 86 3 19 47 65 36 9 38 57 85 
X37 exc-neuron 0 38 67 35 7 33 86 40 69 62 100 65 
X38 exc-neuron 0 39 37 90 68 47 84 27 15 100 53 78 
X39 exc-neuron 0 40 56 26 28 96 69 39 55 73 68 60 
X40 exc-neuron 0 41 66 92 12 28 99 27 36 1 31 32 
X41 exc-neuron 0 42 80 32 17 27 5 54 24 38 51 55 
X42 exc-neuron 0 43 84 35 13 10 73 26 11 6 36 20 
X43 exc-neuron 0 44 65 55 22 47 93 84 27 92 16 9 
X44 exc-neuron 0 45 86 49 8 28 24 89 58 76 2 56 
X45 exc-neuron 0 46 1 72 86 56 34 94 45 16 100 52 
X46 exc-neuron 0 47 44 51 32 43 17 16 41 69 56 63 
X47 exc-neuron 0 48 46 4 68 10 31 9 84 34 93 37 
X48 exc-neuron 0 49 48 7 97 11 61 93 88 74 40 8 
X49 exc-neuron 0 50 3 31 81 25 84 13 39 69 6 78 
X50 exc-neuron 0 51 70 18 81 4 52 82 90 56 19 78 
X51 exc-neuron 0 52 30 26 11 71 8 98 95 32 14 97 
X52 exc-neuron 0 53 82 28 66 92 83 15 72 80 7 30 
X53 exc-neuron 0 54 43 39 100 96 83 74 14 31 79 73 
X54 exc-neuron 0 55 89 12 48 37 21 87 28 9 76 71 
X55 exc-neuron 0 56 16 95 71 9 67 49 97 18 53 37 
X56 exc-neuron 0 57 89 61 52 45 6 14 39 22 64 23 
X57 exc-neuron 0 58 94 84 28 13 61 55 88 100 17 11 
X58 exc-neuron 0 59 32 73 81 29 1 89 56 30 47 48 
X59 exc-neuron 0 60 59 19 72 8 97 37 94 27 76 91 
X60 exc-neuron 0 61 45 30 92 70 39 93 79 56 21 87 
X61 exc-neuron 0 62 5 86 95 49 72 81 64 46 44 82 
X62 exc-neuron 0 63 68 12 25 36 50 40 30 4 74 85 
X63 exc-neuron 0 64 88 55 97 32 5 47 19 29 30 9 
X64 exc-neuron 0 65 35 51 96 15 58 29 52 93 90 61 
X65 exc-neuron 0 66 63 74 50 85 90 97 64 53 32 5 
X66 exc-neuron 0 67 23 81 13 72 14 33 64 19 82 3 
X67 exc-neuron 0 68 62 91 78 59 84 23 38 17 2 30 
X68 exc-neuron 0 69 23 36 95 75 28 35 31 15 70 60 
X69 exc-neuron 0 70 72 32 71 79 53 98 6 44 76 84 
X70 exc-neuron 0 71 81 30 43 80 93 9 66 31 65 13 
X71 exc-neuron 0 72 32 49 93 89 43 38 28 97 51 65 
X72 exc-neuron 0 73 56 99 46 14 13 17 32 21 83 60 
X73 exc-neuron 0 74 47 96 95 42 29 53 60 83 45 23 
X74 exc-neuron 0 75 12 25 69 51 34 48 37 62 6 66 
X75 exc-neuron 0 76 94 44 91 67 40 25 22 63 85 81 
X76 exc-neuron 0 77 68 25 10 50 71 19 53 56 26 40 
X77 exc-neuron 0 78 69 93 76 61 30 68 26 23 40 21 
X78 exc-neuron 0 79 95 56 48 90 34 23 88 49 13 83 
X79 exc-neuron 0 80 66 97 67 47 40 20 56 69 55 65 
X80 exc-neuron 0 81 41 97 84 9 56 61 14 33 95 11 
X81 exc-neuron 0 82 42 27 74 19 29 6 75 67 28 39 
X82 exc-neuron 0 83 41 85 39 59 94 78 93 99 74 37 
X83 exc-neuron 0 84 52 35 51 89 63 8 78 41 61 67 
X84 exc-neuron 0 85 70 25 10 59 88 83 37 34 47 92 
X85 exc-neuron 0 86 22 45 73 5 66 11 17 61 79 59 
X86 exc-neuron 0 87 81 68 33 40 51 32 89 99 92 93 
X87 exc-neuron 0 88 25 43 92 67 77 62 3 4 89 84 
X88 exc-neuron 0 89 86 78 98 62 27 26 74 84 25 68 
X89 exc-neuron 0 90 17 37 94 32 72 16 14 8 10 25 
X90 exc-neuron 0 91 7 30 69 65 29 51 37 85 11 31 
X91 exc-neuron 0 92 93 41 20 70 49 8 86 68 51 87 
X92 exc-neuron 0 93 2 6 61 21 55 79 52 31 56 51 
X93 exc-neuron 0 94 77 33 99 20 16 53 83 37 35 73 
X94 exc-neuron 0 95 73 94 2 15 77 65 48 5 58 93 
X95 exc-neuron 0 96 68 40 25 87 50 60 67 54 73 83 
X96 exc-neuron 0 97 26 4 22 12 3 71 79 80 83 84 
X97 exc-neuron 0 98 22 1 39 44 72 25 64 65 34 70 
X98 exc-neuron 0 99 55 50 3 19 28 21 77 13 89 30 
X99 exc-neuron 0 100 71 46 84 58 59 34 50 19 41 90 

*circuit output 
.tran 0.001p 1049.999p 0 0.001p
.print PHASE B2.X0.X0
.print PHASE B2.X0.X1
.print PHASE B2.X0.X2
.print PHASE B2.X0.X3
.print PHASE B2.X0.X4
.print PHASE B2.X0.X5
.print PHASE B2.X0.X6
.print PHASE B2.X0.X7
.print PHASE B2.X0.X8
.print PHASE B2.X0.X9
.print PHASE B2.X0.X10
.print PHASE B2.X0.X11
.print PHASE B2.X0.X12
.print PHASE B2.X0.X13
.print PHASE B2.X0.X14
.print PHASE B2.X0.X15
.print PHASE B2.X0.X16
.print PHASE B2.X0.X17
.print PHASE B2.X0.X18
.print PHASE B2.X0.X19
.print PHASE B2.X0.X20
.print PHASE B2.X0.X21
.print PHASE B2.X0.X22
.print PHASE B2.X0.X23
.print PHASE B2.X0.X24
.print PHASE B2.X0.X25
.print PHASE B2.X0.X26
.print PHASE B2.X0.X27
.print PHASE B2.X0.X28
.print PHASE B2.X0.X29
.print PHASE B2.X0.X30
.print PHASE B2.X0.X31
.print PHASE B2.X0.X32
.print PHASE B2.X0.X33
.print PHASE B2.X0.X34
.print PHASE B2.X0.X35
.print PHASE B2.X0.X36
.print PHASE B2.X0.X37
.print PHASE B2.X0.X38
.print PHASE B2.X0.X39
.print PHASE B2.X0.X40
.print PHASE B2.X0.X41
.print PHASE B2.X0.X42
.print PHASE B2.X0.X43
.print PHASE B2.X0.X44
.print PHASE B2.X0.X45
.print PHASE B2.X0.X46
.print PHASE B2.X0.X47
.print PHASE B2.X0.X48
.print PHASE B2.X0.X49
.print PHASE B2.X0.X50
.print PHASE B2.X0.X51
.print PHASE B2.X0.X52
.print PHASE B2.X0.X53
.print PHASE B2.X0.X54
.print PHASE B2.X0.X55
.print PHASE B2.X0.X56
.print PHASE B2.X0.X57
.print PHASE B2.X0.X58
.print PHASE B2.X0.X59
.print PHASE B2.X0.X60
.print PHASE B2.X0.X61
.print PHASE B2.X0.X62
.print PHASE B2.X0.X63
.print PHASE B2.X0.X64
.print PHASE B2.X0.X65
.print PHASE B2.X0.X66
.print PHASE B2.X0.X67
.print PHASE B2.X0.X68
.print PHASE B2.X0.X69
.print PHASE B2.X0.X70
.print PHASE B2.X0.X71
.print PHASE B2.X0.X72
.print PHASE B2.X0.X73
.print PHASE B2.X0.X74
.print PHASE B2.X0.X75
.print PHASE B2.X0.X76
.print PHASE B2.X0.X77
.print PHASE B2.X0.X78
.print PHASE B2.X0.X79
.print PHASE B2.X0.X80
.print PHASE B2.X0.X81
.print PHASE B2.X0.X82
.print PHASE B2.X0.X83
.print PHASE B2.X0.X84
.print PHASE B2.X0.X85
.print PHASE B2.X0.X86
.print PHASE B2.X0.X87
.print PHASE B2.X0.X88
.print PHASE B2.X0.X89
.print PHASE B2.X0.X90
.print PHASE B2.X0.X91
.print PHASE B2.X0.X92
.print PHASE B2.X0.X93
.print PHASE B2.X0.X94
.print PHASE B2.X0.X95
.print PHASE B2.X0.X96
.print PHASE B2.X0.X97
.print PHASE B2.X0.X98
.print PHASE B2.X0.X99
.ends
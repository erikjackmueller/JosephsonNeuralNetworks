* Josim Circuit automatically assembled using build_circuit on 2025-09-25 10:36:50.036506 
 
.SUBCKT Neuron-Soma0	0	1	6
* inductances
L0	0	1	3.34pH
L1	2	3	0.51pH
L2	3	4	1.09pH
L3	4	5	4.41pH
L4	5	6	2.21pH

* junctions
B0	1	2	jsoma
B1	4	0	jsoma	
B2	5	0	jsoma ic=250uA

* sources
IB0	0	3	277uA
IB1	0	5	175uA

.model jsoma jj(rtype=0, icrit=225.000uA cap=1.2PF RN=0.925)
.ends Neuron-Soma0

.SUBCKT R-Synapse-exc1	0	1	2
* inductances
R1	1	0	1
RSCALE	1	2	20
.ends R-Synapse-exc1


* main circuit
IIN1 0 1 pwl(0 0 1.892p 0 1.893p 1000000.0u 1.894p 0 2.222p 0 2.223p 1000000.0u 2.224p 0 4.538p 0 4.539p 1000000.0u 4.54p 0 6.764p 0 6.765p 1000000.0u 6.766p 0 8.087p 0 8.088p 1000000.0u 8.089p 0 8.75p 0 8.751p 1000000.0u 8.752p 0 10.028p 0 10.029p 1000000.0u 10.03p 0 11.237p 0 11.238p 1000000.0u 11.239p 0 12.605p 0 12.606p 1000000.0u 12.607p 0 12.77p 0 12.771p 1000000.0u 12.772p 0 17.453p 0 17.454p 1000000.0u 17.455p 0 21.326p 0 21.327p 1000000.0u 21.328p 0 21.83p 0 21.831p 1000000.0u 21.832p 0 29.066p 0 29.067p 1000000.0u 29.068p 0 29.198p 0 29.199p 1000000.0u 29.2p 0 32.171p 0 32.172p 1000000.0u 32.173p 0 35.405p 0 35.406p 1000000.0u 35.407p 0 36.179p 0 36.18p 1000000.0u 36.181p 0 36.299p 0 36.3p 1000000.0u 36.301p 0 37.295p 0 37.296p 1000000.0u 37.297p 0 39.887p 0 39.888p 1000000.0u 39.889p 0 45.869p 0 45.87p 1000000.0u 45.871p 0 46.892p 0 46.893p 1000000.0u 46.894p 0 47.066p 0 47.067p 1000000.0u 47.068p 0 48.323p 0 48.324p 1000000.0u 48.325p 0 53.816p 0 53.817p 1000000.0u 53.818p 0 59.462p 0 59.463p 1000000.0u 59.464p 0 63.524p 0 63.525p 1000000.0u 63.526p 0 63.866p 0 63.867p 1000000.0u 63.868p 0 64.832p 0 64.833p 1000000.0u 64.834p 0 68.567p 0 68.568p 1000000.0u 68.569p 0 70.853p 0 70.854p 1000000.0u 70.855p 0 71.759p 0 71.76p 1000000.0u 71.761p 0 73.979p 0 73.98p 1000000.0u 73.981p 0 75.638p 0 75.639p 1000000.0u 75.64p 0 76.832p 0 76.833p 1000000.0u 76.834p 0 77.948p 0 77.949p 1000000.0u 77.95p 0 78.098p 0 78.099p 1000000.0u 78.1p 0 78.767p 0 78.768p 1000000.0u 78.769p 0 80.621p 0 80.622p 1000000.0u 80.623p 0 80.732p 0 80.733p 1000000.0u 80.734p 0 82.031p 0 82.032p 1000000.0u 82.033p 0 85.187p 0 85.188p 1000000.0u 85.189p 0 85.964p 0 85.965p 1000000.0u 85.966p 0 90.668p 0 90.669p 1000000.0u 90.67p 0 91.394p 0 91.395p 1000000.0u 91.396p 0 93.815p 0 93.816p 1000000.0u 93.817p 0 100.424p 0 100.425p 1000000.0u 100.426p 0 101.753p 0 101.754p 1000000.0u 101.755p 0 106.037p 0 106.038p 1000000.0u 106.039p 0 106.823p 0 106.824p 1000000.0u 106.825p 0 107.702p 0 107.703p 1000000.0u 107.704p 0 108.014p 0 108.015p 1000000.0u 108.016p 0 108.098p 0 108.099p 1000000.0u 108.1p 0 110.294p 0 110.295p 1000000.0u 110.296p 0 111.383p 0 111.384p 1000000.0u 111.385p 0 112.811p 0 112.812p 1000000.0u 112.813p 0 121.667p 0 121.668p 1000000.0u 121.669p 0 126.32p 0 126.321p 1000000.0u 126.322p 0 128.15p 0 128.151p 1000000.0u 128.152p 0 128.84p 0 128.841p 1000000.0u 128.842p 0 129.044p 0 129.045p 1000000.0u 129.046p 0 129.182p 0 129.183p 1000000.0u 129.184p 0 129.923p 0 129.924p 1000000.0u 129.925p 0 130.133p 0 130.134p 1000000.0u 130.135p 0 132.98p 0 132.981p 1000000.0u 132.982p 0 134.333p 0 134.334p 1000000.0u 134.335p 0 137.468p 0 137.469p 1000000.0u 137.47p 0 141.758p 0 141.759p 1000000.0u 141.76p 0 146.39p 0 146.391p 1000000.0u 146.392p 0 149.36p 0 149.361p 1000000.0u 149.362p 0 150.314p 0 150.315p 1000000.0u 150.316p 0 150.626p 0 150.627p 1000000.0u 150.628p 0 151.988p 0 151.989p 1000000.0u 151.99p 0 154.214p 0 154.215p 1000000.0u 154.216p 0 154.994p 0 154.995p 1000000.0u 154.996p 0 155.0p 0 155.001p 1000000.0u 155.002p 0 164.183p 0 164.184p 1000000.0u 164.185p 0 165.95p 0 165.951p 1000000.0u 165.952p 0 166.046p 0 166.047p 1000000.0u 166.048p 0 166.643p 0 166.644p 1000000.0u 166.645p 0 168.794p 0 168.795p 1000000.0u 168.796p 0 168.938p 0 168.939p 1000000.0u 168.94p 0 172.265p 0 172.266p 1000000.0u 172.267p 0 172.328p 0 172.329p 1000000.0u 172.33p 0 174.191p 0 174.192p 1000000.0u 174.193p 0 175.13p 0 175.131p 1000000.0u 175.132p 0 175.433p 0 175.434p 1000000.0u 175.435p 0 178.085p 0 178.086p 1000000.0u 178.087p 0 179.537p 0 179.538p 1000000.0u 179.539p 0 180.221p 0 180.222p 1000000.0u 180.223p 0 181.256p 0 181.257p 1000000.0u 181.258p 0 189.581p 0 189.582p 1000000.0u 189.583p 0 190.091p 0 190.092p 1000000.0u 190.093p 0 190.124p 0 190.125p 1000000.0u 190.126p 0 190.328p 0 190.329p 1000000.0u 190.33p 0 190.358p 0 190.359p 1000000.0u 190.36p 0 191.513p 0 191.514p 1000000.0u 191.515p 0 193.487p 0 193.488p 1000000.0u 193.489p 0 194.714p 0 194.715p 1000000.0u 194.716p 0 195.863p 0 195.864p 1000000.0u 195.865p 0 196.553p 0 196.554p 1000000.0u 196.555p 0 197.771p 0 197.772p 1000000.0u 197.773p 0 199.478p 0 199.479p 1000000.0u 199.48p 0 200.222p 0 200.223p 1000000.0u 200.224p 0 200.669p 0 200.67p 1000000.0u 200.671p 0 201.683p 0 201.684p 1000000.0u 201.685p 0 206.261p 0 206.262p 1000000.0u 206.263p 0 207.791p 0 207.792p 1000000.0u 207.793p 0 211.154p 0 211.155p 1000000.0u 211.156p 0 215.042p 0 215.043p 1000000.0u 215.044p 0 217.937p 0 217.938p 1000000.0u 217.939p 0 219.329p 0 219.33p 1000000.0u 219.331p 0 222.572p 0 222.573p 1000000.0u 222.574p 0 225.182p 0 225.183p 1000000.0u 225.184p 0 225.965p 0 225.966p 1000000.0u 225.967p 0 227.348p 0 227.349p 1000000.0u 227.35p 0 227.549p 0 227.55p 1000000.0u 227.551p 0 227.933p 0 227.934p 1000000.0u 227.935p 0 230.174p 0 230.175p 1000000.0u 230.176p 0 230.639p 0 230.64p 1000000.0u 230.641p 0 235.547p 0 235.548p 1000000.0u 235.549p 0 235.688p 0 235.689p 1000000.0u 235.69p 0 238.901p 0 238.902p 1000000.0u 238.903p 0 239.624p 0 239.625p 1000000.0u 239.626p 0 240.257p 0 240.258p 1000000.0u 240.259p 0 240.263p 0 240.264p 1000000.0u 240.265p 0 242.984p 0 242.985p 1000000.0u 242.986p 0 243.605p 0 243.606p 1000000.0u 243.607p 0 245.537p 0 245.538p 1000000.0u 245.539p 0 246.677p 0 246.678p 1000000.0u 246.679p 0 248.225p 0 248.226p 1000000.0u 248.227p 0 249.656p 0 249.657p 1000000.0u 249.658p 0 251.828p 0 251.829p 1000000.0u 251.83p 0 251.837p 0 251.838p 1000000.0u 251.839p 0 256.736p 0 256.737p 1000000.0u 256.738p 0 256.772p 0 256.773p 1000000.0u 256.774p 0 258.593p 0 258.594p 1000000.0u 258.595p 0 259.043p 0 259.044p 1000000.0u 259.045p 0 260.618p 0 260.619p 1000000.0u 260.62p 0 263.252p 0 263.253p 1000000.0u 263.254p 0 264.374p 0 264.375p 1000000.0u 264.376p 0 264.998p 0 264.999p 1000000.0u 265.0p 0 265.019p 0 265.02p 1000000.0u 265.021p 0 266.471p 0 266.472p 1000000.0u 266.473p 0 266.585p 0 266.586p 1000000.0u 266.587p 0 266.963p 0 266.964p 1000000.0u 266.965p 0 267.248p 0 267.249p 1000000.0u 267.25p 0 268.496p 0 268.497p 1000000.0u 268.498p 0 270.368p 0 270.369p 1000000.0u 270.37p 0 272.006p 0 272.007p 1000000.0u 272.008p 0 273.287p 0 273.288p 1000000.0u 273.289p 0 274.175p 0 274.176p 1000000.0u 274.177p 0 277.472p 0 277.473p 1000000.0u 277.474p 0 279.518p 0 279.519p 1000000.0u 279.52p 0 280.271p 0 280.272p 1000000.0u 280.273p 0 282.308p 0 282.309p 1000000.0u 282.31p 0 283.235p 0 283.236p 1000000.0u 283.237p 0 283.373p 0 283.374p 1000000.0u 283.375p 0 284.483p 0 284.484p 1000000.0u 284.485p 0 284.696p 0 284.697p 1000000.0u 284.698p 0 286.292p 0 286.293p 1000000.0u 286.294p 0 289.232p 0 289.233p 1000000.0u 289.234p 0 292.439p 0 292.44p 1000000.0u 292.441p 0 293.09p 0 293.091p 1000000.0u 293.092p 0 293.114p 0 293.115p 1000000.0u 293.116p 0 294.074p 0 294.075p 1000000.0u 294.076p 0 294.104p 0 294.105p 1000000.0u 294.106p 0 295.133p 0 295.134p 1000000.0u 295.135p 0 297.392p 0 297.393p 1000000.0u 297.394p 0 297.632p 0 297.633p 1000000.0u 297.634p 0 298.085p 0 298.086p 1000000.0u 298.087p 0)

X0 Neuron-Soma0 0 1 2 
X1 R-Synapse-exc1 0 2 3 
ROUT 3 0 1

*circuit output 
.tran 0.001p 319.999p 0 0.001p
.print DEVI IIN1
.print PHASE B0.X0
.print PHASE B1.X0
.print DEVV B0.X0
.print DEVV B1.X0
.print DEVI ROUT
.ends